
module sqroot_comb_NBITS16_DW01_inc_4 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   n1, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n21, n24, n25, n28, n29, n33;

  XOR20 U47 ( .A(n8), .B(n9), .Q(SUM[6]) );
  XOR20 U48 ( .A(n13), .B(n14), .Q(SUM[5]) );
  XOR21 U49 ( .A(n28), .B(n29), .Q(SUM[2]) );
  NAND20 U50 ( .A(A[0]), .B(A[1]), .Q(n29) );
  NAND20 U51 ( .A(A[0]), .B(n25), .Q(n24) );
  NAND20 U52 ( .A(A[0]), .B(n7), .Q(n6) );
  INV2 U53 ( .A(n3), .Q(n2) );
  NOR21 U54 ( .A(n16), .B(n19), .Q(n15) );
  NAND20 U55 ( .A(A[0]), .B(n15), .Q(n14) );
  NAND20 U56 ( .A(A[0]), .B(n10), .Q(n9) );
  INV0 U57 ( .A(n11), .Q(n10) );
  INV2 U58 ( .A(n1), .Q(SUM[8]) );
  INV0 U59 ( .A(n18), .Q(n19) );
  INV0 U60 ( .A(A[5]), .Q(n13) );
  NAND20 U61 ( .A(n7), .B(A[7]), .Q(n3) );
  CLKIN1 U62 ( .A(A[1]), .Q(n33) );
  XOR20 U63 ( .A(n16), .B(n17), .Q(SUM[4]) );
  NOR21 U64 ( .A(n8), .B(n11), .Q(n7) );
  NAND22 U65 ( .A(n18), .B(n12), .Q(n11) );
  NOR21 U66 ( .A(n13), .B(n16), .Q(n12) );
  NOR21 U67 ( .A(n21), .B(n33), .Q(n18) );
  NAND20 U68 ( .A(A[2]), .B(A[3]), .Q(n21) );
  NOR21 U69 ( .A(n28), .B(n33), .Q(n25) );
  INV0 U70 ( .A(A[2]), .Q(n28) );
  INV0 U71 ( .A(A[6]), .Q(n8) );
  NAND20 U72 ( .A(A[0]), .B(n2), .Q(n1) );
  NAND20 U73 ( .A(A[0]), .B(n18), .Q(n17) );
  XNR20 U74 ( .A(A[3]), .B(n24), .Q(SUM[3]) );
  XNR20 U75 ( .A(A[7]), .B(n6), .Q(SUM[7]) );
  INV0 U76 ( .A(A[4]), .Q(n16) );
  XNR20 U77 ( .A(n33), .B(A[0]), .Q(SUM[1]) );
endmodule


module sqroot_comb_NBITS16 ( arg, roundup, sqroot );
  input [15:0] arg;
  output [8:0] sqroot;
  input roundup;
  wire   N711, N712, N713, N714, N715, N716, N717, N718, lt_gt_52_A_7_,
         lt_gt_52_A_4_, lt_gt_52_A_3_, lt_gt_52_A_1_, lt_gt_52_A_0_, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1390,
         n1391, SYNOPSYS_UNCONNECTED_1;

  sqroot_comb_NBITS16_DW01_inc_4 add_53 ( .A({n1391, n746, n1390, n806, n783, 
        lt_gt_52_A_3_, n1121, n757, n646}), .SUM({N718, N717, N716, N715, N714, 
        N713, N712, N711, SYNOPSYS_UNCONNECTED_1}) );
  NAND28 U643 ( .A(n987), .B(n986), .Q(n1047) );
  NAND22 U644 ( .A(n801), .B(n756), .Q(n1281) );
  INV3 U645 ( .A(n1273), .Q(n756) );
  NAND32 U646 ( .A(n1097), .B(n1096), .C(n707), .Q(n1193) );
  INV6 U647 ( .A(n1097), .Q(n1050) );
  NAND21 U648 ( .A(n1196), .B(n673), .Q(n625) );
  INV12 U649 ( .A(n1197), .Q(n685) );
  INV15 U650 ( .A(n1221), .Q(n1273) );
  INV12 U651 ( .A(n815), .Q(n816) );
  INV6 U652 ( .A(n1310), .Q(n1374) );
  NAND22 U653 ( .A(lt_gt_52_A_0_), .B(n1260), .Q(n788) );
  NOR32 U654 ( .A(n1299), .B(n628), .C(n629), .Q(n630) );
  CLKIN3 U655 ( .A(lt_gt_52_A_0_), .Q(n628) );
  CLKIN6 U656 ( .A(n1337), .Q(n1294) );
  NOR23 U657 ( .A(n1390), .B(n1260), .Q(n1227) );
  INV6 U658 ( .A(n631), .Q(n632) );
  INV6 U659 ( .A(n897), .Q(n900) );
  INV10 U660 ( .A(n1034), .Q(n1076) );
  NAND26 U661 ( .A(n653), .B(n870), .Q(n1295) );
  NAND24 U662 ( .A(arg[14]), .B(n811), .Q(n870) );
  NAND32 U663 ( .A(n712), .B(n724), .C(n793), .Q(n653) );
  INV15 U664 ( .A(arg[14]), .Q(n793) );
  OAI2112 U665 ( .A(n1215), .B(n1214), .C(n1213), .D(n1249), .Q(n1216) );
  INV10 U666 ( .A(n1048), .Q(n735) );
  INV2 U667 ( .A(n1048), .Q(n1062) );
  NAND26 U668 ( .A(n1100), .B(n639), .Q(n1148) );
  NAND23 U669 ( .A(n1178), .B(n1177), .Q(n1179) );
  NOR22 U670 ( .A(n1233), .B(n1234), .Q(n798) );
  NAND23 U671 ( .A(n1260), .B(n1390), .Q(n1341) );
  CLKIN10 U672 ( .A(n1188), .Q(n1260) );
  NAND24 U673 ( .A(n1241), .B(n1247), .Q(n1225) );
  NAND24 U674 ( .A(n1276), .B(n1241), .Q(n1252) );
  CLKIN6 U675 ( .A(n1241), .Q(n1218) );
  NAND26 U676 ( .A(n783), .B(n1331), .Q(n1241) );
  INV3 U677 ( .A(n1249), .Q(n1223) );
  NAND23 U678 ( .A(n1298), .B(n784), .Q(n1249) );
  INV3 U679 ( .A(n1274), .Q(n786) );
  AOI212 U680 ( .A(n1066), .B(n1065), .C(n999), .Q(n1002) );
  CLKIN8 U681 ( .A(n1004), .Q(n1075) );
  NAND23 U682 ( .A(n1226), .B(n1225), .Q(n1228) );
  NOR23 U683 ( .A(n1219), .B(n1218), .Q(n1230) );
  CLKIN6 U684 ( .A(n1113), .Q(n1136) );
  NOR32 U685 ( .A(n1233), .B(n1234), .C(n1235), .Q(n1236) );
  NAND34 U686 ( .A(n798), .B(n699), .C(n1348), .Q(n1263) );
  INV2 U687 ( .A(n756), .Q(n757) );
  NAND24 U688 ( .A(n638), .B(n711), .Q(n823) );
  INV4 U689 ( .A(n1031), .Q(n1032) );
  INV6 U690 ( .A(n1076), .Q(n717) );
  INV4 U691 ( .A(n1014), .Q(n1011) );
  NAND24 U692 ( .A(n936), .B(n647), .Q(n1007) );
  INV12 U693 ( .A(n667), .Q(n783) );
  NAND24 U694 ( .A(n960), .B(n906), .Q(n951) );
  NAND42 U695 ( .A(n907), .B(n909), .C(n910), .D(n908), .Q(n973) );
  OAI212 U696 ( .A(n929), .B(n891), .C(n819), .Q(n908) );
  NAND34 U697 ( .A(n945), .B(n944), .C(n806), .Q(n934) );
  INV12 U698 ( .A(n989), .Q(n1064) );
  NOR23 U699 ( .A(n632), .B(n1309), .Q(n1292) );
  CLKIN12 U700 ( .A(n1329), .Q(n815) );
  CLKBU4 U701 ( .A(n1201), .Q(n659) );
  NAND32 U702 ( .A(n967), .B(n966), .C(n981), .Q(n968) );
  CLKIN6 U703 ( .A(n956), .Q(n966) );
  NAND28 U704 ( .A(n1361), .B(n1232), .Q(n1235) );
  XNR22 U705 ( .A(n806), .B(n1345), .Q(n1265) );
  INV3 U706 ( .A(n1201), .Q(n1119) );
  NAND21 U707 ( .A(n1062), .B(n1061), .Q(n626) );
  NAND21 U708 ( .A(n1062), .B(n1061), .Q(n627) );
  NAND28 U709 ( .A(n735), .B(n1061), .Q(n1324) );
  NAND26 U710 ( .A(n1062), .B(n1061), .Q(n1079) );
  BUF2 U711 ( .A(n1079), .Q(n719) );
  CLKIN15 U712 ( .A(n1324), .Q(n1388) );
  CLKIN15 U713 ( .A(n1079), .Q(n1121) );
  NAND28 U714 ( .A(arg[15]), .B(arg[14]), .Q(n820) );
  INV10 U715 ( .A(n678), .Q(n1134) );
  INV6 U716 ( .A(n937), .Q(n1009) );
  NAND34 U717 ( .A(n869), .B(n802), .C(n866), .Q(n944) );
  CLKIN4 U718 ( .A(n869), .Q(n960) );
  CLKIN4 U719 ( .A(n753), .Q(n754) );
  IMUX24 U720 ( .A(n768), .B(n1181), .S(n1273), .Q(n1188) );
  INV6 U721 ( .A(n878), .Q(n894) );
  INV10 U722 ( .A(n1129), .Q(n1186) );
  INV3 U723 ( .A(n1193), .Q(n1204) );
  INV6 U724 ( .A(n944), .Q(n930) );
  NAND22 U725 ( .A(n928), .B(n1355), .Q(n1012) );
  NAND24 U726 ( .A(n696), .B(n850), .Q(n861) );
  NAND22 U727 ( .A(n705), .B(n1089), .Q(n1139) );
  NAND24 U728 ( .A(n876), .B(n879), .Q(n880) );
  BUF12 U729 ( .A(n917), .Q(n802) );
  INV6 U730 ( .A(n916), .Q(n920) );
  NAND23 U731 ( .A(n1091), .B(n1141), .Q(n1088) );
  NOR23 U732 ( .A(n1208), .B(n1209), .Q(n1210) );
  NAND23 U733 ( .A(n1057), .B(n1058), .Q(n1059) );
  NAND22 U734 ( .A(n930), .B(n872), .Q(n648) );
  NAND22 U735 ( .A(n892), .B(n891), .Q(n750) );
  INV3 U736 ( .A(n660), .Q(n751) );
  AOI221 U737 ( .A(arg[15]), .B(arg[12]), .C(n711), .D(n657), .Q(n656) );
  NAND24 U738 ( .A(n847), .B(arg[15]), .Q(n821) );
  NAND33 U739 ( .A(n1070), .B(n782), .C(n1134), .Q(n1102) );
  INV3 U740 ( .A(n1152), .Q(n641) );
  NAND22 U741 ( .A(n930), .B(n693), .Q(n1014) );
  NAND23 U742 ( .A(n1091), .B(n1092), .Q(n1167) );
  NAND22 U743 ( .A(n1072), .B(n1071), .Q(n1078) );
  INV3 U744 ( .A(n803), .Q(n805) );
  INV3 U745 ( .A(n856), .Q(n875) );
  INV3 U746 ( .A(n861), .Q(n853) );
  INV12 U747 ( .A(arg[15]), .Q(n811) );
  NAND24 U748 ( .A(n1358), .B(n1355), .Q(n1361) );
  INV3 U749 ( .A(n1182), .Q(n1340) );
  NAND23 U750 ( .A(n1188), .B(n819), .Q(n1182) );
  INV3 U751 ( .A(n783), .Q(n784) );
  BUF6 U752 ( .A(lt_gt_52_A_7_), .Q(n817) );
  NAND24 U753 ( .A(n1269), .B(n691), .Q(n1296) );
  NOR21 U754 ( .A(n813), .B(n1346), .Q(n1353) );
  INV3 U755 ( .A(n729), .Q(n730) );
  INV3 U756 ( .A(n1041), .Q(n1028) );
  NAND26 U757 ( .A(n1296), .B(n819), .Q(n1297) );
  INV12 U758 ( .A(arg[10]), .Q(n876) );
  INV4 U759 ( .A(n1076), .Q(n651) );
  INV12 U760 ( .A(n804), .Q(lt_gt_52_A_3_) );
  INV12 U761 ( .A(arg[15]), .Q(n810) );
  NOR21 U762 ( .A(n630), .B(n1301), .Q(n1308) );
  INV3 U763 ( .A(n1302), .Q(n629) );
  OAI221 U764 ( .A(lt_gt_52_A_0_), .B(n1300), .C(n1302), .D(n1300), .Q(n1301)
         );
  NOR23 U765 ( .A(n784), .B(n1328), .Q(n631) );
  XNR22 U766 ( .A(n677), .B(n1289), .Q(n1328) );
  NAND22 U767 ( .A(n804), .B(n1286), .Q(n634) );
  NAND22 U768 ( .A(lt_gt_52_A_3_), .B(n633), .Q(n635) );
  NAND22 U769 ( .A(n634), .B(n635), .Q(n1288) );
  INV3 U770 ( .A(n1286), .Q(n633) );
  NAND26 U771 ( .A(lt_gt_52_A_0_), .B(n1288), .Q(n1289) );
  NAND24 U772 ( .A(n636), .B(n637), .Q(n638) );
  CLKIN6 U773 ( .A(arg[11]), .Q(n636) );
  CLKIN6 U774 ( .A(arg[10]), .Q(n637) );
  INV6 U775 ( .A(arg[12]), .Q(n711) );
  BUF6 U776 ( .A(n954), .Q(n721) );
  INV6 U777 ( .A(n706), .Q(n808) );
  NAND23 U778 ( .A(lt_gt_52_A_0_), .B(n1302), .Q(n1279) );
  NAND26 U779 ( .A(n715), .B(n714), .Q(n799) );
  NAND24 U780 ( .A(n1094), .B(n1047), .Q(n1041) );
  NAND24 U781 ( .A(n1184), .B(n783), .Q(n1149) );
  INV6 U782 ( .A(n917), .Q(n919) );
  NAND22 U783 ( .A(n1168), .B(n685), .Q(n1158) );
  INV12 U784 ( .A(n1209), .Q(n1196) );
  INV3 U785 ( .A(n716), .Q(n975) );
  CLKIN1 U786 ( .A(n1213), .Q(n1224) );
  INV6 U787 ( .A(n1261), .Q(n1357) );
  INV8 U788 ( .A(n1264), .Q(n1345) );
  BUF2 U789 ( .A(n678), .Q(n702) );
  NAND26 U790 ( .A(n765), .B(arg[9]), .Q(n917) );
  INV12 U791 ( .A(n1291), .Q(lt_gt_52_A_4_) );
  INV12 U792 ( .A(n683), .Q(n684) );
  NAND24 U793 ( .A(n829), .B(n843), .Q(n834) );
  OAI222 U794 ( .A(n790), .B(n880), .C(n826), .D(n879), .Q(n883) );
  INV15 U795 ( .A(n826), .Q(n790) );
  BUF12 U796 ( .A(n1206), .Q(n639) );
  NAND26 U797 ( .A(n942), .B(n803), .Q(n964) );
  INV10 U798 ( .A(n1122), .Q(n763) );
  INV8 U799 ( .A(n782), .Q(n1141) );
  NOR23 U800 ( .A(n626), .B(n737), .Q(n1084) );
  NAND24 U801 ( .A(n1108), .B(n1109), .Q(n1110) );
  NAND24 U802 ( .A(n898), .B(n640), .Q(n759) );
  CLKBU12 U803 ( .A(n826), .Q(n652) );
  INV12 U804 ( .A(arg[13]), .Q(n710) );
  IMUX22 U805 ( .A(n774), .B(n1063), .S(n1388), .Q(n1133) );
  CLKIN6 U806 ( .A(n1156), .Q(n1168) );
  NAND24 U807 ( .A(n733), .B(n1153), .Q(n1156) );
  INV6 U808 ( .A(n1347), .Q(n1359) );
  NAND26 U809 ( .A(n1263), .B(n1262), .Q(n1329) );
  CLKIN6 U810 ( .A(n982), .Q(n1015) );
  NAND34 U811 ( .A(n1041), .B(n1042), .C(lt_gt_52_A_3_), .Q(n1043) );
  NAND22 U812 ( .A(n664), .B(n1336), .Q(n1058) );
  NAND28 U813 ( .A(n868), .B(n694), .Q(n862) );
  INV4 U814 ( .A(n851), .Q(n655) );
  NAND33 U815 ( .A(n651), .B(n668), .C(n1053), .Q(n1021) );
  INV6 U816 ( .A(n1052), .Q(n1053) );
  NAND26 U817 ( .A(n881), .B(n882), .Q(n658) );
  NAND34 U818 ( .A(n831), .B(n832), .C(arg[10]), .Q(n881) );
  NAND21 U819 ( .A(n894), .B(n819), .Q(n888) );
  NAND26 U820 ( .A(lt_gt_52_A_4_), .B(n904), .Q(n916) );
  INV15 U821 ( .A(n817), .Q(n1355) );
  NAND23 U822 ( .A(n863), .B(n876), .Q(n882) );
  INV12 U823 ( .A(n781), .Q(n782) );
  NAND28 U824 ( .A(n876), .B(n879), .Q(n849) );
  INV15 U825 ( .A(arg[11]), .Q(n879) );
  OAI312 U826 ( .A(n793), .B(n811), .C(n701), .D(n846), .Q(n852) );
  NAND24 U827 ( .A(n712), .B(n710), .Q(n701) );
  NAND24 U828 ( .A(arg[14]), .B(n810), .Q(n857) );
  INV6 U829 ( .A(n676), .Q(n832) );
  IMUX24 U830 ( .A(n679), .B(n680), .S(n1388), .Q(n678) );
  NAND23 U831 ( .A(n695), .B(n656), .Q(n709) );
  INV8 U832 ( .A(n1093), .Q(n1115) );
  OAI211 U833 ( .A(arg[4]), .B(n1093), .C(arg[5]), .Q(n1201) );
  BUF6 U834 ( .A(n800), .Q(n780) );
  OAI310 U835 ( .A(n847), .B(n811), .C(n701), .D(n846), .Q(n642) );
  AOI222 U836 ( .A(arg[12]), .B(arg[13]), .C(arg[13]), .D(n810), .Q(n846) );
  NAND22 U837 ( .A(n944), .B(n927), .Q(n935) );
  NAND33 U838 ( .A(n712), .B(n724), .C(n793), .Q(n871) );
  XNR21 U839 ( .A(n904), .B(n790), .Q(n901) );
  INV3 U840 ( .A(n1030), .Q(n1033) );
  INV6 U841 ( .A(n927), .Q(n872) );
  INV3 U842 ( .A(n1202), .Q(n1212) );
  NOR22 U843 ( .A(arg[13]), .B(arg[12]), .Q(n839) );
  CLKIN6 U844 ( .A(n766), .Q(n767) );
  NAND23 U845 ( .A(n861), .B(n817), .Q(n766) );
  INV12 U846 ( .A(n1329), .Q(lt_gt_52_A_0_) );
  INV6 U847 ( .A(n867), .Q(n893) );
  NAND23 U848 ( .A(n767), .B(n860), .Q(n867) );
  NOR21 U849 ( .A(n658), .B(n819), .Q(n697) );
  INV3 U850 ( .A(n738), .Q(n739) );
  NOR21 U851 ( .A(arg[6]), .B(n1015), .Q(n738) );
  INV3 U852 ( .A(n759), .Q(n760) );
  INV6 U853 ( .A(n1096), .Q(n1051) );
  NAND22 U854 ( .A(n930), .B(n872), .Q(n936) );
  NAND22 U855 ( .A(n904), .B(lt_gt_52_A_4_), .Q(n905) );
  INV3 U856 ( .A(n890), .Q(n770) );
  NAND22 U857 ( .A(n911), .B(n1355), .Q(n909) );
  INV3 U858 ( .A(n1007), .Q(n747) );
  INV6 U859 ( .A(n763), .Q(n674) );
  INV3 U860 ( .A(n700), .Q(n679) );
  NAND23 U861 ( .A(n747), .B(n746), .Q(n748) );
  NAND22 U862 ( .A(n933), .B(n819), .Q(n1008) );
  CLKIN3 U863 ( .A(n935), .Q(n933) );
  CLKIN12 U864 ( .A(n779), .Q(n991) );
  INV3 U865 ( .A(n703), .Q(n913) );
  INV3 U866 ( .A(n909), .Q(n914) );
  INV3 U867 ( .A(n852), .Q(n695) );
  INV3 U868 ( .A(n849), .Q(n657) );
  INV3 U869 ( .A(n884), .Q(n843) );
  NAND24 U870 ( .A(n712), .B(n724), .Q(n848) );
  IMUX22 U871 ( .A(n1212), .B(n1211), .S(n1210), .Q(n1298) );
  INV3 U872 ( .A(n692), .Q(n693) );
  NAND24 U873 ( .A(lt_gt_52_A_3_), .B(n1290), .Q(n1276) );
  INV3 U874 ( .A(n1000), .Q(n990) );
  XNR21 U875 ( .A(arg[4]), .B(n1121), .Q(n1199) );
  INV3 U876 ( .A(n1046), .Q(n672) );
  AOI211 U877 ( .A(n1045), .B(n805), .C(n1044), .Q(n1046) );
  INV3 U878 ( .A(n1150), .Q(n1127) );
  NAND22 U879 ( .A(n1122), .B(n1336), .Q(n1150) );
  NAND23 U880 ( .A(n743), .B(n742), .Q(n745) );
  NAND22 U881 ( .A(n655), .B(n695), .Q(n696) );
  NAND23 U882 ( .A(n708), .B(n709), .Q(n850) );
  NAND22 U883 ( .A(n642), .B(n704), .Q(n708) );
  INV12 U884 ( .A(arg[14]), .Q(n847) );
  NAND22 U885 ( .A(n1355), .B(n761), .Q(n705) );
  INV3 U886 ( .A(n1157), .Q(n1163) );
  NAND26 U887 ( .A(n767), .B(n661), .Q(n694) );
  NAND26 U888 ( .A(n825), .B(n794), .Q(n840) );
  NAND23 U889 ( .A(n811), .B(n793), .Q(n794) );
  NAND22 U890 ( .A(n847), .B(n810), .Q(lt_gt_52_A_7_) );
  CLKIN6 U891 ( .A(n1253), .Q(n1266) );
  NAND24 U892 ( .A(n726), .B(n1336), .Q(n1333) );
  XNR21 U893 ( .A(n1312), .B(n801), .Q(n1325) );
  INV6 U894 ( .A(n1372), .Q(n1375) );
  NOR22 U895 ( .A(n1368), .B(n1369), .Q(n729) );
  BUF6 U896 ( .A(n652), .Q(n806) );
  INV15 U897 ( .A(n903), .Q(n891) );
  NAND22 U898 ( .A(n934), .B(n721), .Q(n938) );
  INV3 U899 ( .A(n1064), .Q(n668) );
  BUF12 U900 ( .A(n921), .Q(n758) );
  CLKIN6 U901 ( .A(n1065), .Q(n1056) );
  OAI222 U902 ( .A(n784), .B(n734), .C(n1175), .D(n1174), .Q(n1178) );
  NAND24 U903 ( .A(n998), .B(n652), .Q(n1054) );
  INV3 U904 ( .A(n1154), .Q(n732) );
  INV3 U905 ( .A(n1263), .Q(n1254) );
  INV6 U906 ( .A(n1164), .Q(n1159) );
  INV6 U907 ( .A(n1200), .Q(n1118) );
  NAND24 U908 ( .A(n1259), .B(n789), .Q(n1261) );
  INV2 U909 ( .A(n1067), .Q(n998) );
  AOI222 U910 ( .A(n963), .B(n964), .C(n1064), .D(n1295), .Q(n962) );
  NOR33 U911 ( .A(n1081), .B(n1080), .C(n627), .Q(n1082) );
  NAND24 U912 ( .A(n1294), .B(n1293), .Q(n1384) );
  INV3 U913 ( .A(n628), .Q(n646) );
  NAND22 U914 ( .A(n964), .B(n963), .Q(n1006) );
  INV6 U915 ( .A(n1295), .Q(n1390) );
  INV3 U916 ( .A(n1314), .Q(lt_gt_52_A_1_) );
  INV3 U917 ( .A(n1339), .Q(n690) );
  INV3 U918 ( .A(n1047), .Q(n996) );
  INV3 U919 ( .A(n1177), .Q(n1155) );
  CLKBU12 U920 ( .A(n1127), .Q(n762) );
  INV6 U921 ( .A(n1213), .Q(n1247) );
  XOR22 U922 ( .A(n819), .B(n658), .Q(n640) );
  INV6 U923 ( .A(n891), .Q(n749) );
  INV3 U924 ( .A(n1095), .Q(n707) );
  AOI211 U925 ( .A(n1255), .B(n1390), .C(n1254), .Q(n1257) );
  INV6 U926 ( .A(n1148), .Q(n1175) );
  NAND22 U927 ( .A(n1365), .B(n798), .Q(n1380) );
  INV3 U928 ( .A(n1172), .Q(n1070) );
  NAND21 U929 ( .A(n1253), .B(n1336), .Q(n1339) );
  INV4 U930 ( .A(n763), .Q(n755) );
  NAND28 U931 ( .A(n655), .B(n787), .Q(n826) );
  CLKIN0 U932 ( .A(n1043), .Q(n1044) );
  CLKIN6 U933 ( .A(n1090), .Q(n1151) );
  INV6 U934 ( .A(n1298), .Q(n1331) );
  INV6 U935 ( .A(n1258), .Q(n1255) );
  INV3 U936 ( .A(n1088), .Q(n1103) );
  NAND22 U937 ( .A(n1167), .B(n819), .Q(n1157) );
  INV6 U938 ( .A(n1107), .Q(n1108) );
  OAI212 U939 ( .A(n992), .B(n991), .C(n1052), .Q(n664) );
  NAND26 U940 ( .A(n992), .B(n991), .Q(n1052) );
  NAND24 U941 ( .A(n713), .B(n891), .Q(n715) );
  INV0 U942 ( .A(n1331), .Q(n740) );
  NAND21 U943 ( .A(n1102), .B(n1136), .Q(n1140) );
  XOR31 U944 ( .A(n664), .B(n727), .C(n1068), .Q(n680) );
  INV12 U945 ( .A(n806), .Q(n1336) );
  NAND28 U946 ( .A(n1196), .B(n673), .Q(n1197) );
  NAND22 U947 ( .A(arg[8]), .B(lt_gt_52_A_4_), .Q(n918) );
  INV0 U948 ( .A(n951), .Q(n952) );
  OAI211 U949 ( .A(n884), .B(n883), .C(n658), .Q(n887) );
  NAND23 U950 ( .A(n1315), .B(n1314), .Q(n1318) );
  INV12 U951 ( .A(n1207), .Q(n1208) );
  BUF2 U952 ( .A(n1306), .Q(n643) );
  NOR33 U953 ( .A(n1319), .B(n1121), .C(n816), .Q(n1320) );
  INV1 U954 ( .A(n1345), .Q(n807) );
  IMUX22 U955 ( .A(n723), .B(n1360), .S(n1359), .Q(n1362) );
  NAND21 U956 ( .A(n1258), .B(n819), .Q(n1256) );
  XOR22 U957 ( .A(n666), .B(n746), .Q(n1346) );
  CLKIN2 U958 ( .A(n1380), .Q(n1367) );
  NAND24 U959 ( .A(n815), .B(n1304), .Q(n1305) );
  OAI212 U960 ( .A(arg[0]), .B(n682), .C(arg[1]), .Q(n1317) );
  AOI212 U961 ( .A(n1364), .B(n1363), .C(n1362), .Q(n1365) );
  XNR22 U962 ( .A(n741), .B(n1279), .Q(n644) );
  NOR23 U963 ( .A(n1291), .B(n770), .Q(n769) );
  NOR22 U964 ( .A(n1291), .B(n770), .Q(n654) );
  CLKBU4 U965 ( .A(n1283), .Q(n645) );
  NAND24 U966 ( .A(n1187), .B(n719), .Q(n1283) );
  INV2 U967 ( .A(n1379), .Q(n665) );
  INV12 U968 ( .A(n991), .Q(n1069) );
  INV0 U969 ( .A(n950), .Q(n953) );
  CLKIN2 U970 ( .A(n930), .Q(n669) );
  OAI2112 U971 ( .A(arg[11]), .B(n652), .C(n658), .D(n1355), .Q(n885) );
  NAND21 U972 ( .A(n1281), .B(n1282), .Q(n1303) );
  NAND24 U973 ( .A(n1043), .B(n997), .Q(n1065) );
  NAND22 U974 ( .A(n945), .B(n669), .Q(n946) );
  INV10 U975 ( .A(n967), .Q(n957) );
  NOR23 U976 ( .A(n730), .B(n1370), .Q(n1371) );
  AOI312 U977 ( .A(n1377), .B(n665), .C(n1367), .D(n1366), .Q(n1368) );
  NOR24 U978 ( .A(n764), .B(n842), .Q(n844) );
  INV6 U979 ( .A(n1297), .Q(n1309) );
  INV1 U980 ( .A(n970), .Q(n994) );
  XOR31 U981 ( .A(n1390), .B(n1167), .C(n1156), .Q(n1169) );
  NAND21 U982 ( .A(n659), .B(n812), .Q(n1202) );
  INV3 U983 ( .A(n943), .Q(n647) );
  INV3 U984 ( .A(n928), .Q(n943) );
  NAND22 U985 ( .A(n899), .B(n900), .Q(n928) );
  NOR23 U986 ( .A(n1069), .B(n1064), .Q(n649) );
  XOR22 U987 ( .A(n769), .B(n780), .Q(n650) );
  NAND24 U988 ( .A(n905), .B(n802), .Q(n949) );
  OAI211 U989 ( .A(n1028), .B(n1040), .C(n1027), .Q(n1029) );
  NAND28 U990 ( .A(n877), .B(n827), .Q(n828) );
  NAND28 U991 ( .A(n831), .B(n832), .Q(n877) );
  OAI222 U992 ( .A(n848), .B(n821), .C(n820), .D(n710), .Q(n851) );
  NAND23 U993 ( .A(n958), .B(n959), .Q(n778) );
  INV15 U994 ( .A(n1208), .Q(n673) );
  NAND23 U995 ( .A(n881), .B(n882), .Q(n833) );
  NAND24 U996 ( .A(n841), .B(n840), .Q(n787) );
  NAND20 U997 ( .A(n658), .B(n819), .Q(n895) );
  CLKIN15 U998 ( .A(n803), .Q(n804) );
  INV8 U999 ( .A(n1287), .Q(n803) );
  AOI212 U1000 ( .A(n841), .B(n840), .C(n851), .Q(n842) );
  NAND28 U1001 ( .A(n840), .B(n841), .Q(n831) );
  NOR21 U1002 ( .A(n1314), .B(n1272), .Q(n1214) );
  XOR21 U1003 ( .A(n757), .B(n1313), .Q(n1319) );
  INV2 U1004 ( .A(n1387), .Q(sqroot[8]) );
  NOR24 U1005 ( .A(n892), .B(n891), .Q(n660) );
  INV6 U1006 ( .A(n929), .Q(n892) );
  INV4 U1007 ( .A(n958), .Q(n776) );
  NOR24 U1008 ( .A(n957), .B(n718), .Q(n958) );
  IMUX23 U1009 ( .A(n875), .B(n874), .S(n790), .Q(n661) );
  IMUX23 U1010 ( .A(n875), .B(n874), .S(n790), .Q(n860) );
  INV6 U1011 ( .A(n828), .Q(n835) );
  NAND24 U1012 ( .A(n1113), .B(n1112), .Q(n1207) );
  CLKIN4 U1013 ( .A(n844), .Q(n743) );
  XNR22 U1014 ( .A(n892), .B(n749), .Q(n931) );
  INV2 U1015 ( .A(n1242), .Q(n1243) );
  BUF2 U1016 ( .A(n796), .Q(n662) );
  NOR21 U1017 ( .A(n668), .B(n1053), .Q(n663) );
  CLKIN6 U1018 ( .A(n668), .Q(n774) );
  OAI211 U1019 ( .A(n992), .B(n991), .C(n1052), .Q(n1067) );
  INV3 U1020 ( .A(n1102), .Q(n1104) );
  NAND23 U1021 ( .A(n763), .B(n806), .Q(n1128) );
  OAI211 U1022 ( .A(n1364), .B(n1363), .C(n1354), .Q(n1377) );
  INV6 U1023 ( .A(n1376), .Q(n1379) );
  CLKIN2 U1024 ( .A(n1359), .Q(n666) );
  CLKIN4 U1025 ( .A(lt_gt_52_A_4_), .Q(n667) );
  NAND21 U1026 ( .A(n955), .B(n721), .Q(n959) );
  NAND34 U1027 ( .A(n799), .B(n1012), .C(n1390), .Q(n978) );
  NAND21 U1028 ( .A(n1076), .B(n1324), .Q(n1077) );
  NOR24 U1029 ( .A(n697), .B(n893), .Q(n896) );
  NAND42 U1030 ( .A(n1114), .B(n1096), .C(n707), .D(n1097), .Q(n706) );
  XOR22 U1031 ( .A(n677), .B(n1289), .Q(n670) );
  INV3 U1032 ( .A(n785), .Q(n677) );
  XOR22 U1033 ( .A(n1255), .B(n1390), .Q(n1259) );
  INV1 U1034 ( .A(n1223), .Q(n671) );
  CLKIN2 U1035 ( .A(n1184), .Q(n734) );
  NAND23 U1036 ( .A(n996), .B(n995), .Q(n1042) );
  NAND20 U1037 ( .A(n1042), .B(n1041), .Q(n1045) );
  INV6 U1038 ( .A(n1101), .Q(n1203) );
  OAI222 U1039 ( .A(n675), .B(n981), .C(n980), .D(n716), .Q(n983) );
  MUX26 U1040 ( .A(n996), .B(n672), .S(n1115), .Q(n1129) );
  INV2 U1041 ( .A(n650), .Q(n675) );
  NAND34 U1042 ( .A(n951), .B(n950), .C(n783), .Q(n954) );
  INV6 U1043 ( .A(n966), .Q(n718) );
  OAI222 U1044 ( .A(n848), .B(n821), .C(n820), .D(n710), .Q(n676) );
  NAND22 U1045 ( .A(n681), .B(n1173), .Q(n1154) );
  NAND20 U1046 ( .A(n801), .B(n719), .Q(n1321) );
  NAND24 U1047 ( .A(n1061), .B(n735), .Q(n773) );
  NAND32 U1048 ( .A(n1091), .B(n1092), .C(n1390), .Q(n1164) );
  NAND34 U1049 ( .A(n1196), .B(n1272), .C(n673), .Q(n1242) );
  NAND24 U1050 ( .A(n644), .B(n727), .Q(n728) );
  CLKIN6 U1051 ( .A(n1231), .Q(n1358) );
  NAND28 U1052 ( .A(n823), .B(n684), .Q(n841) );
  INV6 U1053 ( .A(n762), .Q(n681) );
  NAND22 U1054 ( .A(n877), .B(n876), .Q(n878) );
  OAI222 U1055 ( .A(arg[6]), .B(n995), .C(n805), .D(n981), .Q(n969) );
  NAND22 U1056 ( .A(arg[6]), .B(n978), .Q(n980) );
  CLKIN2 U1057 ( .A(lt_gt_52_A_0_), .Q(n682) );
  NAND23 U1058 ( .A(n1172), .B(n702), .Q(n1092) );
  INV15 U1059 ( .A(arg[13]), .Q(n724) );
  NAND23 U1060 ( .A(n1036), .B(n1035), .Q(n1048) );
  NAND26 U1061 ( .A(n868), .B(n694), .Q(n1291) );
  NAND23 U1062 ( .A(n869), .B(n866), .Q(n950) );
  NAND24 U1063 ( .A(lt_gt_52_A_3_), .B(n1327), .Q(n1307) );
  NOR22 U1064 ( .A(n1280), .B(n804), .Q(n1219) );
  CLKIN6 U1065 ( .A(n1086), .Q(n1091) );
  OAI211 U1066 ( .A(lt_gt_52_A_1_), .B(n1272), .C(n1282), .Q(n1277) );
  NAND20 U1067 ( .A(n973), .B(n978), .Q(n977) );
  INV3 U1068 ( .A(n1175), .Q(n731) );
  NAND28 U1069 ( .A(n822), .B(n824), .Q(n683) );
  NAND24 U1070 ( .A(n1198), .B(n685), .Q(n686) );
  NAND23 U1071 ( .A(n1197), .B(n1199), .Q(n687) );
  NAND26 U1072 ( .A(n686), .B(n687), .Q(n688) );
  CLKIN12 U1073 ( .A(n688), .Q(n1280) );
  NAND22 U1074 ( .A(n689), .B(n690), .Q(n691) );
  INV0 U1075 ( .A(n1345), .Q(n689) );
  INV12 U1076 ( .A(n862), .Q(n902) );
  INV2 U1077 ( .A(n918), .Q(n915) );
  NAND24 U1078 ( .A(n931), .B(n943), .Q(n692) );
  OAI211 U1079 ( .A(n953), .B(n952), .C(n784), .Q(n955) );
  NAND22 U1080 ( .A(n994), .B(n784), .Q(n1066) );
  INV1 U1081 ( .A(n1232), .Q(n698) );
  INV2 U1082 ( .A(n698), .Q(n699) );
  INV6 U1083 ( .A(n795), .Q(n1232) );
  NAND32 U1084 ( .A(n1171), .B(n1172), .C(n806), .Q(n1090) );
  INV6 U1085 ( .A(n1176), .Q(n1184) );
  INV0 U1086 ( .A(n1006), .Q(n1022) );
  BUF2 U1087 ( .A(n1069), .Q(n700) );
  INV6 U1088 ( .A(n1087), .Q(n1160) );
  OAI2110 U1089 ( .A(n1022), .B(n1021), .C(lt_gt_52_A_3_), .D(n1020), .Q(n1023) );
  NAND20 U1090 ( .A(n1022), .B(n1021), .Q(n1144) );
  INV2 U1091 ( .A(n639), .Q(n1194) );
  OAI212 U1092 ( .A(n919), .B(n920), .C(n1336), .Q(n703) );
  OAI222 U1093 ( .A(n811), .B(n711), .C(arg[12]), .D(n849), .Q(n704) );
  NAND21 U1094 ( .A(n1064), .B(n819), .Q(n775) );
  NAND28 U1095 ( .A(n900), .B(n899), .Q(n911) );
  NAND28 U1096 ( .A(n902), .B(n760), .Q(n899) );
  NAND32 U1097 ( .A(n868), .B(n694), .C(n865), .Q(n765) );
  OAI222 U1098 ( .A(n774), .B(n1053), .C(n649), .D(n1052), .Q(n1060) );
  NOR20 U1099 ( .A(n1222), .B(n625), .Q(n1220) );
  INV6 U1100 ( .A(n921), .Q(n922) );
  BUF2 U1101 ( .A(n960), .Q(n720) );
  INV6 U1102 ( .A(n968), .Q(n993) );
  NAND23 U1103 ( .A(n844), .B(n845), .Q(n744) );
  NAND22 U1104 ( .A(n831), .B(arg[11]), .Q(n829) );
  NAND26 U1105 ( .A(n871), .B(n870), .Q(n884) );
  NOR33 U1106 ( .A(n739), .B(n975), .C(n985), .Q(n976) );
  OAI2112 U1107 ( .A(n1028), .B(n1040), .C(n783), .D(n1027), .Q(n997) );
  INV8 U1108 ( .A(n864), .Q(n868) );
  INV15 U1109 ( .A(arg[12]), .Q(n712) );
  NAND22 U1110 ( .A(n903), .B(n892), .Q(n714) );
  INV2 U1111 ( .A(n892), .Q(n713) );
  IMUX24 U1112 ( .A(n752), .B(n1185), .S(n1273), .Q(n1253) );
  OAI212 U1113 ( .A(n914), .B(n913), .C(n758), .Q(n716) );
  NAND26 U1114 ( .A(n777), .B(n778), .Q(n779) );
  INV3 U1115 ( .A(n1098), .Q(n1099) );
  NAND24 U1116 ( .A(n912), .B(n818), .Q(n921) );
  INV6 U1117 ( .A(n911), .Q(n912) );
  NAND21 U1118 ( .A(n1013), .B(n1012), .Q(n1016) );
  INV1 U1119 ( .A(n980), .Q(n984) );
  IMUX24 U1120 ( .A(n722), .B(n1169), .S(n1273), .Q(n1231) );
  BUF2 U1121 ( .A(n702), .Q(n722) );
  BUF2 U1122 ( .A(n1361), .Q(n723) );
  NAND24 U1123 ( .A(n1088), .B(n1102), .Q(n1087) );
  NAND24 U1124 ( .A(n950), .B(n949), .Q(n945) );
  INV2 U1125 ( .A(n974), .Q(n985) );
  XOR22 U1126 ( .A(n1355), .B(n1075), .Q(n737) );
  NAND22 U1127 ( .A(n725), .B(lt_gt_52_A_0_), .Q(n726) );
  CLKIN2 U1128 ( .A(n1330), .Q(n725) );
  NAND24 U1129 ( .A(n728), .B(n1335), .Q(n1372) );
  INV1 U1130 ( .A(n1336), .Q(n727) );
  XOR22 U1131 ( .A(n814), .B(n1333), .Q(n1334) );
  INV2 U1132 ( .A(n1381), .Q(n1369) );
  XNR22 U1133 ( .A(n646), .B(n1371), .Q(sqroot[0]) );
  NAND33 U1134 ( .A(n1177), .B(n731), .C(n732), .Q(n733) );
  NOR33 U1135 ( .A(n1355), .B(n1104), .C(n1103), .Q(n1105) );
  NAND33 U1136 ( .A(n735), .B(n1061), .C(n1124), .Q(n1097) );
  NAND21 U1137 ( .A(n1171), .B(n1172), .Q(n1180) );
  BUF2 U1138 ( .A(n1348), .Q(n736) );
  INV3 U1139 ( .A(n1170), .Q(n1348) );
  NAND21 U1140 ( .A(n935), .B(n648), .Q(n873) );
  CLKIN15 U1141 ( .A(n1027), .Q(n992) );
  BUF12 U1142 ( .A(n1295), .Q(n819) );
  XOR22 U1143 ( .A(n1242), .B(n1049), .Q(n1187) );
  NOR22 U1144 ( .A(n1329), .B(n1265), .Q(n1267) );
  CLKIN1 U1145 ( .A(n755), .Q(n768) );
  NAND24 U1146 ( .A(n748), .B(n932), .Q(n941) );
  INV3 U1147 ( .A(n740), .Q(n741) );
  NAND24 U1148 ( .A(n745), .B(n744), .Q(n854) );
  INV3 U1149 ( .A(n845), .Q(n742) );
  NAND22 U1150 ( .A(n1066), .B(n1065), .Q(n1068) );
  CLKIN3 U1151 ( .A(n1355), .Q(n746) );
  NAND28 U1152 ( .A(n750), .B(n751), .Q(n927) );
  BUF2 U1153 ( .A(n1186), .Q(n752) );
  INV6 U1154 ( .A(n1283), .Q(n1248) );
  NAND28 U1155 ( .A(n1196), .B(n673), .Q(n1221) );
  NAND33 U1156 ( .A(n935), .B(n648), .C(n1390), .Q(n937) );
  NAND20 U1157 ( .A(n1390), .B(n1000), .Q(n1001) );
  NAND22 U1158 ( .A(n649), .B(n992), .Q(n1000) );
  INV3 U1159 ( .A(n1054), .Q(n999) );
  CLKIN2 U1160 ( .A(n1252), .Q(n753) );
  NAND20 U1161 ( .A(n740), .B(n806), .Q(n1299) );
  INV2 U1162 ( .A(n1118), .Q(n812) );
  INV2 U1163 ( .A(n1276), .Q(n1274) );
  AOI310 U1164 ( .A(n1121), .B(n1222), .C(n1314), .D(n1220), .Q(n1229) );
  XNR22 U1165 ( .A(n783), .B(n1278), .Q(n1330) );
  NAND22 U1166 ( .A(n966), .B(n967), .Q(n1287) );
  NAND20 U1167 ( .A(n1015), .B(n1014), .Q(n1018) );
  NAND26 U1168 ( .A(n1280), .B(n804), .Q(n1213) );
  AOI212 U1169 ( .A(n954), .B(n934), .C(n797), .Q(n796) );
  NAND28 U1170 ( .A(n902), .B(n901), .Q(n903) );
  XNR22 U1171 ( .A(arg[11]), .B(n894), .Q(n898) );
  CLKIN2 U1172 ( .A(n1160), .Q(n761) );
  NAND24 U1173 ( .A(n1121), .B(n1306), .Q(n1285) );
  OAI211 U1174 ( .A(n1355), .B(n1103), .C(n1163), .Q(n1089) );
  NAND24 U1175 ( .A(n876), .B(n884), .Q(n764) );
  AOI212 U1176 ( .A(n1253), .B(n1336), .C(n1223), .Q(n1226) );
  NAND34 U1177 ( .A(n1186), .B(n763), .C(n808), .Q(n1172) );
  NAND24 U1178 ( .A(n775), .B(n965), .Q(n1038) );
  NAND28 U1179 ( .A(n1047), .B(n792), .Q(n1027) );
  NAND34 U1180 ( .A(n974), .B(n979), .C(n982), .Q(n967) );
  NAND24 U1181 ( .A(n1115), .B(n1094), .Q(n1200) );
  XOR22 U1182 ( .A(arg[2]), .B(n685), .Q(n801) );
  NAND22 U1183 ( .A(lt_gt_52_A_0_), .B(n1311), .Q(n1312) );
  XOR22 U1184 ( .A(arg[12]), .B(n857), .Q(n858) );
  NAND28 U1185 ( .A(arg[12]), .B(arg[14]), .Q(n824) );
  NAND28 U1186 ( .A(arg[12]), .B(arg[13]), .Q(n822) );
  INV2 U1187 ( .A(n877), .Q(n837) );
  NAND33 U1188 ( .A(n1034), .B(n1006), .C(n818), .Q(n1035) );
  NOR21 U1189 ( .A(arg[5]), .B(n1095), .Q(n771) );
  NOR33 U1190 ( .A(n772), .B(n1050), .C(n1051), .Q(n1101) );
  INV3 U1191 ( .A(n771), .Q(n772) );
  NAND28 U1192 ( .A(n773), .B(arg[4]), .Q(n1096) );
  NAND24 U1193 ( .A(n720), .B(n776), .Q(n777) );
  NAND23 U1194 ( .A(n1266), .B(n806), .Q(n1240) );
  INV6 U1195 ( .A(n1280), .Q(n1290) );
  AOI212 U1196 ( .A(n1303), .B(n1285), .C(n1284), .Q(n1286) );
  NAND21 U1197 ( .A(n741), .B(n1336), .Q(n1332) );
  OAI210 U1198 ( .A(n707), .B(n1199), .C(n1193), .Q(n1195) );
  CLKIN6 U1199 ( .A(n1133), .Q(n781) );
  NAND22 U1200 ( .A(n812), .B(n659), .Q(n1098) );
  CLKIN6 U1201 ( .A(n1252), .Q(n1246) );
  INV3 U1202 ( .A(n1078), .Q(n1081) );
  NAND21 U1203 ( .A(n1221), .B(n1141), .Q(n1351) );
  AOI2111 U1204 ( .A(n1168), .B(n1164), .C(n1221), .D(n1163), .Q(n1166) );
  NOR42 U1205 ( .A(n1159), .B(n1151), .C(n1106), .D(n1105), .Q(n1107) );
  INV6 U1206 ( .A(n1117), .Q(n1126) );
  OAI211 U1207 ( .A(n1204), .B(n1212), .C(n1203), .Q(n1205) );
  INV10 U1208 ( .A(n1386), .Q(n1385) );
  XNR22 U1209 ( .A(n643), .B(n1305), .Q(n1327) );
  OAI211 U1210 ( .A(n1129), .B(n1203), .C(n674), .Q(n1171) );
  NAND23 U1211 ( .A(n949), .B(n1336), .Q(n939) );
  NOR41 U1212 ( .A(n678), .B(n1203), .C(n1129), .D(n755), .Q(n1086) );
  NOR32 U1213 ( .A(n1118), .B(n1119), .C(n804), .Q(n1120) );
  AOI212 U1214 ( .A(n1121), .B(arg[4]), .C(n1120), .Q(n1123) );
  OAI222 U1215 ( .A(n784), .B(n1129), .C(n1126), .D(n1125), .Q(n1131) );
  CLKIN2 U1216 ( .A(n1072), .Q(n1073) );
  OAI221 U1217 ( .A(n1384), .B(n1338), .C(n1337), .D(n1372), .Q(n1370) );
  INV2 U1218 ( .A(n788), .Q(n789) );
  OAI2112 U1219 ( .A(n1204), .B(n1099), .C(n1203), .D(lt_gt_52_A_3_), .Q(n1100) );
  OAI222 U1220 ( .A(n1390), .B(n1134), .C(n818), .D(n782), .Q(n1135) );
  BUF2 U1221 ( .A(n1290), .Q(n785) );
  AOI312 U1222 ( .A(n1277), .B(n786), .C(n1285), .D(n1275), .Q(n1278) );
  OAI212 U1223 ( .A(n1274), .B(n645), .C(n1213), .Q(n1275) );
  INV2 U1224 ( .A(n939), .Q(n797) );
  INV2 U1225 ( .A(n791), .Q(n792) );
  NOR21 U1226 ( .A(n1074), .B(n1073), .Q(n1085) );
  INV3 U1227 ( .A(arg[7]), .Q(n988) );
  NAND20 U1228 ( .A(n1094), .B(n988), .Q(n791) );
  INV1 U1229 ( .A(n1385), .Q(n809) );
  CLKIN2 U1230 ( .A(n1016), .Q(n1019) );
  CLKIN3 U1231 ( .A(n1332), .Q(n814) );
  OAI210 U1232 ( .A(n662), .B(n1009), .C(n1008), .Q(n1010) );
  AOI210 U1233 ( .A(n690), .B(n1341), .C(n1340), .Q(n1342) );
  CLKIN1 U1234 ( .A(n1071), .Q(n1074) );
  INV3 U1235 ( .A(n1077), .Q(n1083) );
  NAND43 U1236 ( .A(n1147), .B(n1351), .C(n1349), .D(n1350), .Q(n795) );
  XNR31 U1237 ( .A(n1184), .B(n783), .C(n1183), .Q(n1185) );
  OAI310 U1238 ( .A(n1142), .B(n719), .C(n1026), .D(n1025), .Q(n1233) );
  OAI310 U1239 ( .A(n1011), .B(n1355), .C(n747), .D(n1010), .Q(n1013) );
  NAND24 U1240 ( .A(n1162), .B(n1161), .Q(n1349) );
  INV3 U1241 ( .A(n1281), .Q(n1245) );
  BUF2 U1242 ( .A(lt_gt_52_A_7_), .Q(n818) );
  AOI210 U1243 ( .A(n1195), .B(n1079), .C(n1194), .Q(n1198) );
  INV0 U1244 ( .A(n1283), .Q(n1284) );
  MUX21 U1245 ( .A(n875), .B(n874), .S(n790), .Q(n800) );
  NOR20 U1246 ( .A(n1364), .B(n1363), .Q(n1352) );
  NOR21 U1247 ( .A(arg[2]), .B(n1313), .Q(n1215) );
  NOR21 U1248 ( .A(arg[8]), .B(n906), .Q(n907) );
  INV3 U1249 ( .A(n857), .Q(n838) );
  AOI211 U1250 ( .A(arg[11]), .B(n1295), .C(n1355), .Q(n889) );
  LOGIC0 U1251 ( .Q(n1391) );
  AOI2112 U1252 ( .A(n1183), .B(n641), .C(n762), .D(n1155), .Q(n1106) );
  MUX21 U1253 ( .A(N717), .B(n746), .S(n1385), .Q(sqroot[7]) );
  INV2 U1254 ( .A(n1296), .Q(n1270) );
  OAI210 U1255 ( .A(n1355), .B(n1004), .C(n1078), .Q(n1005) );
  OAI212 U1256 ( .A(n1118), .B(n1116), .C(n804), .Q(n1117) );
  INV3 U1257 ( .A(n1330), .Q(n1302) );
  AOI312 U1258 ( .A(n802), .B(n806), .C(n905), .D(n915), .Q(n925) );
  IMUX24 U1259 ( .A(n949), .B(n948), .S(n947), .Q(n989) );
  NOR24 U1260 ( .A(n718), .B(n957), .Q(n947) );
  NAND22 U1261 ( .A(n1188), .B(n1295), .Q(n1189) );
  XNR22 U1262 ( .A(arg[3]), .B(n1243), .Q(n1306) );
  NAND21 U1263 ( .A(n1231), .B(n746), .Q(n1170) );
  XNR22 U1264 ( .A(n780), .B(n654), .Q(n982) );
  NAND30 U1265 ( .A(n1350), .B(n1351), .C(n1349), .Q(n1363) );
  BUF2 U1266 ( .A(n1358), .Q(n813) );
  AOI312 U1267 ( .A(n784), .B(n1128), .C(n1129), .D(n1127), .Q(n1130) );
  XNR22 U1268 ( .A(n1321), .B(n1320), .Q(n1322) );
  NAND21 U1269 ( .A(n1373), .B(n1374), .Q(n1338) );
  NAND22 U1270 ( .A(n1031), .B(n1030), .Q(n971) );
  XNR22 U1271 ( .A(arg[7]), .B(n993), .Q(n1040) );
  XNR22 U1272 ( .A(arg[12]), .B(n827), .Q(n856) );
  INV6 U1273 ( .A(n880), .Q(n827) );
  AOI211 U1274 ( .A(n1115), .B(n1124), .C(n1114), .Q(n1116) );
  IMUX24 U1275 ( .A(n1040), .B(n1039), .S(n1115), .Q(n1122) );
  INV6 U1276 ( .A(n1149), .Q(n1152) );
  XNR22 U1277 ( .A(n865), .B(n862), .Q(n869) );
  XNR22 U1278 ( .A(n941), .B(n940), .Q(n942) );
  IMUX22 U1279 ( .A(n1268), .B(n1267), .S(n1266), .Q(n1269) );
  NAND28 U1280 ( .A(n972), .B(n971), .Q(n1061) );
  NOR33 U1281 ( .A(n1136), .B(n1135), .C(n1137), .Q(n1209) );
  XNR22 U1282 ( .A(arg[7]), .B(n993), .Q(n970) );
  IMUX24 U1283 ( .A(n927), .B(n926), .S(n803), .Q(n1034) );
  XNR22 U1284 ( .A(n1355), .B(n1160), .Q(n1165) );
  MUX21 U1285 ( .A(N711), .B(lt_gt_52_A_1_), .S(n1385), .Q(sqroot[1]) );
  MUX21 U1286 ( .A(N712), .B(n1121), .S(n1385), .Q(sqroot[2]) );
  MUX21 U1287 ( .A(N713), .B(lt_gt_52_A_3_), .S(n1385), .Q(sqroot[3]) );
  MUX21 U1288 ( .A(N714), .B(n783), .S(n1385), .Q(sqroot[4]) );
  MUX21 U1289 ( .A(N715), .B(n806), .S(n1385), .Q(sqroot[5]) );
  MUX21 U1290 ( .A(N716), .B(n1390), .S(n1385), .Q(sqroot[6]) );
  XNR22 U1291 ( .A(n1355), .B(n1075), .Q(n1080) );
  OAI222 U1292 ( .A(n810), .B(n710), .C(arg[13]), .D(arg[15]), .Q(n825) );
  XNR21 U1293 ( .A(arg[10]), .B(n790), .Q(n929) );
  CLKIN3 U1294 ( .A(arg[9]), .Q(n830) );
  CLKIN3 U1295 ( .A(arg[8]), .Q(n865) );
  NAND22 U1296 ( .A(n830), .B(n865), .Q(n863) );
  OAI212 U1297 ( .A(n834), .B(n835), .C(n833), .Q(n836) );
  OAI312 U1298 ( .A(n817), .B(n837), .C(n856), .D(n836), .Q(n855) );
  OAI212 U1299 ( .A(n839), .B(n838), .C(arg[11]), .Q(n845) );
  NOR33 U1300 ( .A(n853), .B(n854), .C(n855), .Q(n864) );
  OAI212 U1301 ( .A(arg[13]), .B(arg[14]), .C(n858), .Q(n859) );
  CLKIN3 U1302 ( .A(n859), .Q(n874) );
  CLKIN3 U1303 ( .A(n863), .Q(n904) );
  CLKIN3 U1304 ( .A(arg[6]), .Q(n981) );
  NAND22 U1305 ( .A(n981), .B(n988), .Q(n906) );
  CLKIN3 U1306 ( .A(n906), .Q(n866) );
  XOR31 U1307 ( .A(n1390), .B(n796), .C(n873), .Q(n926) );
  OAI212 U1308 ( .A(n818), .B(n1390), .C(n885), .Q(n886) );
  AOI312 U1309 ( .A(n889), .B(n888), .C(n887), .D(n886), .Q(n890) );
  OAI222 U1310 ( .A(n896), .B(n898), .C(n895), .D(n898), .Q(n897) );
  OAI212 U1311 ( .A(n919), .B(n920), .C(n1336), .Q(n910) );
  OAI222 U1312 ( .A(n978), .B(n650), .C(n973), .D(n650), .Q(n956) );
  OAI212 U1313 ( .A(n914), .B(n913), .C(n758), .Q(n979) );
  OAI312 U1314 ( .A(n1336), .B(n919), .C(n920), .D(n918), .Q(n923) );
  AOI212 U1315 ( .A(n799), .B(n923), .C(n922), .Q(n924) );
  OAI212 U1316 ( .A(n1295), .B(n925), .C(n924), .Q(n974) );
  AOI212 U1317 ( .A(n1007), .B(n1355), .C(n1011), .Q(n932) );
  AOI312 U1318 ( .A(n939), .B(n1008), .C(n938), .D(n1009), .Q(n940) );
  NAND22 U1319 ( .A(n1287), .B(n943), .Q(n963) );
  XOR31 U1320 ( .A(n1336), .B(n954), .C(n946), .Q(n948) );
  OAI222 U1321 ( .A(n1336), .B(n1069), .C(n1064), .D(n1295), .Q(n961) );
  OAI2112 U1322 ( .A(n818), .B(n1034), .C(n962), .D(n961), .Q(n1036) );
  AOI222 U1323 ( .A(n1069), .B(n1336), .C(n964), .D(n963), .Q(n965) );
  AOI212 U1324 ( .A(n1076), .B(n1355), .C(n1038), .Q(n972) );
  CLKIN3 U1325 ( .A(arg[4]), .Q(n1124) );
  CLKIN3 U1326 ( .A(arg[5]), .Q(n1114) );
  NAND22 U1327 ( .A(n1124), .B(n1114), .Q(n995) );
  OAI212 U1328 ( .A(n970), .B(n783), .C(n969), .Q(n1031) );
  NAND22 U1329 ( .A(n970), .B(n783), .Q(n1030) );
  CLKIN3 U1330 ( .A(n995), .Q(n1094) );
  AOI312 U1331 ( .A(n675), .B(n981), .C(n977), .D(n976), .Q(n987) );
  AOI212 U1332 ( .A(n985), .B(n984), .C(n983), .Q(n986) );
  OAI212 U1333 ( .A(n990), .B(n651), .C(n1021), .Q(n1004) );
  NAND22 U1334 ( .A(n663), .B(n819), .Q(n1071) );
  CLKIN3 U1335 ( .A(n1058), .Q(n1003) );
  OAI222 U1336 ( .A(n1003), .B(n1002), .C(n663), .D(n1001), .Q(n1072) );
  OAI212 U1337 ( .A(n818), .B(n1075), .C(n1005), .Q(n1142) );
  CLKIN3 U1338 ( .A(n1018), .Q(n1017) );
  OAI222 U1339 ( .A(n1019), .B(n1018), .C(n1017), .D(n1016), .Q(n1020) );
  NAND22 U1340 ( .A(n1144), .B(n1023), .Q(n1026) );
  CLKIN3 U1341 ( .A(n1144), .Q(n1143) );
  CLKIN3 U1342 ( .A(n1023), .Q(n1024) );
  OAI212 U1343 ( .A(n1143), .B(n1142), .C(n1024), .Q(n1025) );
  XOR31 U1344 ( .A(n783), .B(n1043), .C(n1029), .Q(n1039) );
  OAI222 U1345 ( .A(n717), .B(n818), .C(n1032), .D(n1033), .Q(n1037) );
  OAI2112 U1346 ( .A(n1038), .B(n1037), .C(n1036), .D(n1035), .Q(n1093) );
  CLKIN3 U1347 ( .A(arg[3]), .Q(n1049) );
  CLKIN3 U1348 ( .A(arg[2]), .Q(n1272) );
  NAND22 U1349 ( .A(n1049), .B(n1272), .Q(n1095) );
  CLKIN3 U1350 ( .A(n1066), .Q(n1055) );
  OAI212 U1351 ( .A(n1056), .B(n1055), .C(n1054), .Q(n1057) );
  XOR31 U1352 ( .A(n1390), .B(n1060), .C(n1059), .Q(n1063) );
  AOI2112 U1353 ( .A(n1085), .B(n1084), .C(n1083), .D(n1082), .Q(n1113) );
  CLKIN3 U1354 ( .A(n1140), .Q(n1109) );
  NAND22 U1355 ( .A(n1098), .B(n804), .Q(n1173) );
  OAI2112 U1356 ( .A(arg[4]), .B(n707), .C(n1193), .D(n1121), .Q(n1206) );
  NAND22 U1357 ( .A(n1173), .B(n1148), .Q(n1183) );
  OAI222 U1358 ( .A(n1186), .B(n808), .C(n1203), .D(n1129), .Q(n1176) );
  NAND22 U1359 ( .A(n1176), .B(n784), .Q(n1177) );
  OAI222 U1360 ( .A(n1139), .B(n1110), .C(n1109), .D(n1108), .Q(n1138) );
  OAI2112 U1361 ( .A(arg[15]), .B(n782), .C(n1390), .D(n1134), .Q(n1111) );
  OAI212 U1362 ( .A(n1355), .B(n1141), .C(n1111), .Q(n1112) );
  OAI222 U1363 ( .A(n1126), .B(n1123), .C(n1336), .D(n674), .Q(n1132) );
  NAND22 U1364 ( .A(n707), .B(n1124), .Q(n1125) );
  OAI212 U1365 ( .A(n1132), .B(n1131), .C(n1130), .Q(n1137) );
  NAND22 U1366 ( .A(n1196), .B(n673), .Q(n1314) );
  AOI2112 U1367 ( .A(n1140), .B(n1139), .C(n1314), .D(n1138), .Q(n1234) );
  CLKIN3 U1368 ( .A(n1142), .Q(n1145) );
  OAI222 U1369 ( .A(n1145), .B(n1144), .C(n1143), .D(n1142), .Q(n1146) );
  NAND22 U1370 ( .A(n1121), .B(n1146), .Q(n1147) );
  CLKIN3 U1371 ( .A(n1147), .Q(n1354) );
  OAI212 U1372 ( .A(n1152), .B(n1151), .C(n681), .Q(n1153) );
  OAI222 U1373 ( .A(n1158), .B(n1159), .C(n1157), .D(n1221), .Q(n1162) );
  CLKIN6 U1374 ( .A(n1165), .Q(n1161) );
  NAND22 U1375 ( .A(n1166), .B(n1165), .Q(n1350) );
  CLKIN3 U1376 ( .A(n1173), .Q(n1174) );
  XOR31 U1377 ( .A(n806), .B(n1180), .C(n1179), .Q(n1181) );
  OAI212 U1378 ( .A(n1340), .B(n1240), .C(n1341), .Q(n1239) );
  AOI212 U1379 ( .A(n1253), .B(n1336), .C(n1248), .Q(n1190) );
  NAND24 U1380 ( .A(n1190), .B(n1189), .Q(n1217) );
  CLKIN3 U1381 ( .A(arg[1]), .Q(n1192) );
  CLKIN3 U1382 ( .A(arg[0]), .Q(n1191) );
  NAND22 U1383 ( .A(n1192), .B(n1191), .Q(n1313) );
  XOR31 U1384 ( .A(n639), .B(lt_gt_52_A_3_), .C(n1205), .Q(n1211) );
  NOR24 U1385 ( .A(n1217), .B(n1216), .Q(n1238) );
  NAND22 U1386 ( .A(arg[3]), .B(n1121), .Q(n1222) );
  AOI2112 U1387 ( .A(n1230), .B(n1229), .C(n1227), .D(n1228), .Q(n1237) );
  OAI312 U1388 ( .A(n1239), .B(n1238), .C(n1237), .D(n1236), .Q(n1262) );
  CLKIN3 U1389 ( .A(n1240), .Q(n1344) );
  NAND22 U1390 ( .A(n1313), .B(n1272), .Q(n1282) );
  CLKIN3 U1391 ( .A(n1282), .Q(n1244) );
  OAI212 U1392 ( .A(n1245), .B(n1244), .C(n1285), .Q(n1251) );
  OAI212 U1393 ( .A(n1248), .B(n1224), .C(n1246), .Q(n1250) );
  OAI2112 U1394 ( .A(n754), .B(n1251), .C(n1250), .D(n671), .Q(n1264) );
  OAI212 U1395 ( .A(n1344), .B(n1345), .C(n1339), .Q(n1258) );
  OAI222 U1396 ( .A(n1260), .B(n1257), .C(n1260), .D(n1256), .Q(n1356) );
  OAI212 U1397 ( .A(n1336), .B(n807), .C(n815), .Q(n1268) );
  CLKIN3 U1398 ( .A(roundup), .Q(n1366) );
  AOI212 U1399 ( .A(n1270), .B(n1390), .C(n1366), .Q(n1271) );
  OAI312 U1400 ( .A(n1356), .B(n1355), .C(n1357), .D(n1271), .Q(n1337) );
  OAI212 U1401 ( .A(n806), .B(n644), .C(n1292), .Q(n1293) );
  NAND22 U1402 ( .A(n1299), .B(n806), .Q(n1300) );
  XNR21 U1403 ( .A(n1303), .B(n1121), .Q(n1304) );
  OAI222 U1404 ( .A(n1309), .B(n1308), .C(n1309), .D(n1307), .Q(n1310) );
  CLKIN3 U1405 ( .A(n1319), .Q(n1311) );
  NAND22 U1406 ( .A(n1329), .B(arg[0]), .Q(n1316) );
  OAI212 U1407 ( .A(n1313), .B(n816), .C(n1316), .Q(n1315) );
  AOI222 U1408 ( .A(n1318), .B(n1317), .C(lt_gt_52_A_1_), .D(n1316), .Q(n1323)
         );
  OAI222 U1409 ( .A(n1325), .B(n719), .C(n1323), .D(n1322), .Q(n1326) );
  OAI2112 U1410 ( .A(lt_gt_52_A_3_), .B(n1327), .C(n1326), .D(n1297), .Q(n1373) );
  OAI212 U1411 ( .A(n783), .B(n670), .C(n1334), .Q(n1335) );
  CLKIN3 U1412 ( .A(n1341), .Q(n1343) );
  OAI312 U1413 ( .A(n1343), .B(n1344), .C(n1345), .D(n1342), .Q(n1347) );
  OAI212 U1414 ( .A(n736), .B(n1359), .C(n723), .Q(n1364) );
  OAI2112 U1415 ( .A(n1353), .B(n1352), .C(n646), .D(roundup), .Q(n1381) );
  OAI212 U1416 ( .A(n1357), .B(n1356), .C(n1355), .Q(n1376) );
  NAND22 U1417 ( .A(n813), .B(n746), .Q(n1360) );
  OAI222 U1418 ( .A(n1375), .B(n1374), .C(n1373), .D(n1375), .Q(n1383) );
  CLKIN3 U1419 ( .A(n1377), .Q(n1378) );
  OAI312 U1420 ( .A(n1380), .B(n1379), .C(n1378), .D(roundup), .Q(n1382) );
  OAI2112 U1421 ( .A(n1384), .B(n1383), .C(n1382), .D(n1381), .Q(n1386) );
  NAND22 U1422 ( .A(N718), .B(n809), .Q(n1387) );
endmodule

