
module sqroot_comb_NBITS32_DW01_sub_28 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n3, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n33, n34, n35, n38, n40, n43, n45, n47, n48, n49, n50,
         n51, n53, n54, n55, n56, n58, n59, n60, n62, n63, n65, n66, n67, n70,
         n72, n75, n77, n79, n82, n83, n86, n88, n91, n92, n93, n95, n96, n99,
         n101, n104, n108, n110, n113, n116, n118, n121, n123, n125, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n145, n146, n147, n148, n149, n150, n151, n152, n155,
         n156, n157, n158, n159, n161, n162, n163, n164, n165, n166, n167,
         n168, n171, n172, n173, n174, n175, n176, n177, n180, n181, n182,
         n183, n184, n185, n186, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n210,
         n211, n212, n213, n214, n215, n218, n219, n220, n222, n223, n224,
         n225, n226, n228, n229, n230, n231, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n246, n247, n254, n257, n259, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405;

  OAI212 U38 ( .A(n393), .B(n391), .C(n58), .Q(n56) );
  OAI212 U63 ( .A(n394), .B(n391), .C(n77), .Q(n75) );
  OAI212 U83 ( .A(n394), .B(n391), .C(n93), .Q(n91) );
  OAI212 U121 ( .A(n394), .B(n391), .C(n123), .Q(n121) );
  OAI212 U155 ( .A(n147), .B(n196), .C(n148), .Q(n146) );
  OAI212 U163 ( .A(n163), .B(n155), .C(n156), .Q(n150) );
  OAI212 U179 ( .A(n364), .B(n196), .C(n370), .Q(n164) );
  AOI212 U185 ( .A(n171), .B(n186), .C(n172), .Q(n166) );
  OAI212 U203 ( .A(n183), .B(n196), .C(n184), .Q(n182) );
  NAND28 U295 ( .A(n375), .B(n374), .Q(n376) );
  AOI211 U296 ( .A(n225), .B(n246), .C(n222), .Q(n220) );
  NOR21 U297 ( .A(A[21]), .B(A[20]), .Q(n96) );
  OAI211 U298 ( .A(n394), .B(n391), .C(n101), .Q(n99) );
  XNR21 U299 ( .A(n20), .B(n157), .Q(DIFF[14]) );
  NAND23 U300 ( .A(n185), .B(n171), .Q(n165) );
  CLKIN4 U301 ( .A(n391), .Q(n381) );
  NAND21 U302 ( .A(n391), .B(n384), .Q(n382) );
  INV12 U303 ( .A(n197), .Q(n196) );
  INV2 U304 ( .A(n186), .Q(n184) );
  AOI211 U305 ( .A(n168), .B(n238), .C(n161), .Q(n159) );
  NOR23 U306 ( .A(n165), .B(n131), .Q(n129) );
  BUF2 U307 ( .A(n374), .Q(n362) );
  NAND20 U308 ( .A(n239), .B(n174), .Q(n22) );
  NAND24 U309 ( .A(n388), .B(n174), .Q(n172) );
  INV4 U310 ( .A(n150), .Q(n152) );
  NOR24 U311 ( .A(n404), .B(A[4]), .Q(n229) );
  OAI211 U312 ( .A(n394), .B(n391), .C(n53), .Q(n51) );
  CLKIN2 U313 ( .A(n184), .Q(n367) );
  INV8 U314 ( .A(n226), .Q(n225) );
  INV2 U315 ( .A(n152), .Q(n366) );
  NAND22 U316 ( .A(n242), .B(n195), .Q(n25) );
  NAND24 U317 ( .A(A[9]), .B(n396), .Q(n195) );
  NAND26 U318 ( .A(n149), .B(n133), .Q(n131) );
  INV1 U319 ( .A(A[26]), .Q(n62) );
  NOR23 U320 ( .A(n108), .B(n82), .Q(n77) );
  INV4 U321 ( .A(n142), .Q(n236) );
  CLKIN6 U322 ( .A(n236), .Q(n365) );
  NOR24 U323 ( .A(n397), .B(A[13]), .Q(n162) );
  NAND24 U324 ( .A(n225), .B(n385), .Q(n386) );
  AOI211 U325 ( .A(n367), .B(n240), .C(n387), .Q(n177) );
  INV6 U326 ( .A(n374), .Q(n379) );
  INV6 U327 ( .A(n230), .Q(n228) );
  CLKIN6 U328 ( .A(n229), .Q(n247) );
  XNR21 U329 ( .A(A[31]), .B(n31), .Q(DIFF[31]) );
  INV3 U330 ( .A(n19), .Q(n380) );
  INV3 U331 ( .A(n21), .Q(n373) );
  XNR21 U332 ( .A(A[30]), .B(n38), .Q(DIFF[30]) );
  NAND22 U333 ( .A(n236), .B(n145), .Q(n19) );
  INV3 U334 ( .A(n167), .Q(n364) );
  NAND21 U335 ( .A(n392), .B(n123), .Q(n17) );
  INV0 U336 ( .A(n123), .Q(n125) );
  XOR21 U337 ( .A(n211), .B(n27), .Q(DIFF[7]) );
  NAND21 U338 ( .A(n60), .B(n55), .Q(n54) );
  CLKIN3 U339 ( .A(n392), .Q(n393) );
  NAND23 U340 ( .A(n48), .B(n77), .Q(n47) );
  NOR24 U341 ( .A(n401), .B(A[16]), .Q(n377) );
  NAND21 U342 ( .A(A[14]), .B(n398), .Q(n156) );
  NOR21 U343 ( .A(A[18]), .B(A[19]), .Q(n113) );
  OAI212 U344 ( .A(n365), .B(n152), .C(n145), .Q(n141) );
  CLKIN0 U345 ( .A(n194), .Q(n242) );
  NAND23 U346 ( .A(A[17]), .B(n402), .Q(n123) );
  NAND22 U347 ( .A(n167), .B(n149), .Q(n147) );
  INV3 U348 ( .A(n149), .Q(n151) );
  CLKIN3 U349 ( .A(n191), .Q(n241) );
  NAND22 U350 ( .A(A[6]), .B(n259), .Q(n219) );
  NOR23 U351 ( .A(n191), .B(n194), .Q(n185) );
  INV3 U352 ( .A(n92), .Q(n392) );
  INV1 U353 ( .A(n185), .Q(n183) );
  BUF2 U354 ( .A(n213), .Q(n363) );
  INV6 U355 ( .A(n165), .Q(n167) );
  AOI212 U356 ( .A(n200), .B(n213), .C(n201), .Q(n199) );
  NAND23 U357 ( .A(A[15]), .B(n395), .Q(n145) );
  XNR21 U358 ( .A(A[28]), .B(n51), .Q(DIFF[28]) );
  NAND21 U359 ( .A(n50), .B(n55), .Q(n49) );
  NAND20 U360 ( .A(n362), .B(n219), .Q(n28) );
  NAND24 U361 ( .A(A[11]), .B(n254), .Q(n181) );
  INV2 U362 ( .A(n180), .Q(n240) );
  INV1 U363 ( .A(n214), .Q(n368) );
  CLKIN3 U364 ( .A(n212), .Q(n214) );
  INV4 U365 ( .A(n207), .Q(n244) );
  INV6 U366 ( .A(n381), .Q(n369) );
  INV2 U367 ( .A(n168), .Q(n370) );
  INV6 U368 ( .A(n166), .Q(n168) );
  NAND26 U369 ( .A(A[7]), .B(n403), .Q(n210) );
  NAND22 U370 ( .A(A[8]), .B(n257), .Q(n203) );
  CLKIN4 U371 ( .A(n244), .Q(n371) );
  OAI211 U372 ( .A(n371), .B(n215), .C(n210), .Q(n206) );
  XNR22 U373 ( .A(A[25]), .B(n70), .Q(DIFF[25]) );
  INV2 U374 ( .A(n213), .Q(n215) );
  NOR23 U375 ( .A(n254), .B(A[11]), .Q(n180) );
  CLKIN12 U376 ( .A(n218), .Q(n374) );
  NOR24 U377 ( .A(n259), .B(A[6]), .Q(n218) );
  XNR21 U378 ( .A(A[29]), .B(n43), .Q(DIFF[29]) );
  NAND24 U379 ( .A(n67), .B(n62), .Q(n59) );
  INV1 U380 ( .A(n223), .Q(n246) );
  NAND22 U381 ( .A(A[16]), .B(n401), .Q(n136) );
  NAND23 U382 ( .A(A[4]), .B(n404), .Q(n230) );
  NAND24 U383 ( .A(n387), .B(n239), .Q(n388) );
  CLKIN6 U384 ( .A(n198), .Q(n385) );
  NAND24 U385 ( .A(n212), .B(n200), .Q(n198) );
  NAND21 U386 ( .A(n240), .B(n181), .Q(n23) );
  OAI211 U387 ( .A(n394), .B(n391), .C(n65), .Q(n63) );
  NAND28 U388 ( .A(A[5]), .B(n405), .Q(n224) );
  AOI212 U389 ( .A(n168), .B(n149), .C(n366), .Q(n148) );
  CLKIN12 U390 ( .A(n224), .Q(n375) );
  INV0 U391 ( .A(n202), .Q(n243) );
  INV6 U392 ( .A(n181), .Q(n387) );
  NOR21 U393 ( .A(n371), .B(n214), .Q(n205) );
  XNR21 U394 ( .A(A[24]), .B(n75), .Q(DIFF[24]) );
  CLKIN3 U395 ( .A(B[9]), .Q(n396) );
  NAND24 U396 ( .A(n113), .B(n123), .Q(n108) );
  NOR21 U397 ( .A(n54), .B(n79), .Q(n53) );
  CLKIN6 U398 ( .A(n77), .Q(n79) );
  INV10 U399 ( .A(n197), .Q(n372) );
  XOR22 U400 ( .A(n164), .B(n373), .Q(DIFF[13]) );
  XNR22 U401 ( .A(A[19]), .B(n116), .Q(DIFF[19]) );
  NAND22 U402 ( .A(A[10]), .B(n399), .Q(n192) );
  NOR24 U403 ( .A(n399), .B(A[10]), .Q(n191) );
  OAI211 U404 ( .A(n393), .B(n369), .C(n33), .Q(n31) );
  OAI211 U405 ( .A(n394), .B(n369), .C(n40), .Q(n38) );
  NAND28 U406 ( .A(n376), .B(n219), .Q(n213) );
  XOR22 U407 ( .A(n28), .B(n220), .Q(DIFF[6]) );
  NAND21 U408 ( .A(n243), .B(n203), .Q(n26) );
  INV6 U409 ( .A(n173), .Q(n239) );
  INV1 U410 ( .A(n47), .Q(n45) );
  INV1 U411 ( .A(A[27]), .Q(n55) );
  OAI211 U412 ( .A(n393), .B(n391), .C(n45), .Q(n43) );
  NOR23 U413 ( .A(n405), .B(A[5]), .Q(n223) );
  NAND22 U414 ( .A(A[12]), .B(n400), .Q(n174) );
  CLKBU15 U415 ( .A(n2), .Q(n391) );
  NOR21 U416 ( .A(A[24]), .B(A[25]), .Q(n67) );
  XOR20 U417 ( .A(n372), .B(n25), .Q(DIFF[9]) );
  NAND20 U418 ( .A(A[5]), .B(n405), .Q(n378) );
  NOR24 U419 ( .A(n162), .B(n155), .Q(n149) );
  XOR22 U420 ( .A(n380), .B(n146), .Q(DIFF[15]) );
  NAND21 U421 ( .A(n237), .B(n156), .Q(n20) );
  OAI212 U422 ( .A(n393), .B(n391), .C(n118), .Q(n116) );
  XNR22 U423 ( .A(n23), .B(n182), .Q(DIFF[11]) );
  NOR24 U424 ( .A(n400), .B(A[12]), .Q(n173) );
  OAI212 U425 ( .A(n194), .B(n372), .C(n195), .Q(n193) );
  OAI212 U426 ( .A(n138), .B(n372), .C(n139), .Q(n137) );
  NAND21 U427 ( .A(n167), .B(n140), .Q(n138) );
  NOR24 U428 ( .A(n202), .B(n207), .Q(n200) );
  NOR24 U429 ( .A(n403), .B(A[7]), .Q(n207) );
  NOR22 U430 ( .A(n396), .B(A[9]), .Q(n194) );
  NAND24 U431 ( .A(n381), .B(n17), .Q(n383) );
  NAND24 U432 ( .A(n382), .B(n383), .Q(DIFF[17]) );
  INV3 U433 ( .A(n17), .Q(n384) );
  AOI212 U434 ( .A(n150), .B(n133), .C(n134), .Q(n132) );
  NOR24 U435 ( .A(n377), .B(n142), .Q(n133) );
  XNR21 U436 ( .A(A[21]), .B(n99), .Q(DIFF[21]) );
  NAND21 U437 ( .A(n235), .B(n136), .Q(n18) );
  XNR22 U438 ( .A(A[23]), .B(n86), .Q(DIFF[23]) );
  NOR21 U439 ( .A(n59), .B(n79), .Q(n58) );
  NAND28 U440 ( .A(n386), .B(n199), .Q(n197) );
  NOR24 U441 ( .A(n257), .B(A[8]), .Q(n202) );
  INV2 U442 ( .A(n378), .Q(n222) );
  NAND21 U443 ( .A(n246), .B(n378), .Q(n29) );
  XNR22 U444 ( .A(n22), .B(n175), .Q(DIFF[12]) );
  OAI212 U445 ( .A(n393), .B(n391), .C(n72), .Q(n70) );
  NOR22 U446 ( .A(n365), .B(n151), .Q(n140) );
  OAI212 U447 ( .A(n145), .B(n135), .C(n136), .Q(n134) );
  XNR22 U448 ( .A(n24), .B(n193), .Q(DIFF[10]) );
  XNR22 U449 ( .A(n18), .B(n137), .Q(DIFF[16]) );
  NOR23 U450 ( .A(n173), .B(n180), .Q(n171) );
  XNR22 U451 ( .A(n121), .B(A[18]), .Q(DIFF[18]) );
  NOR21 U452 ( .A(n402), .B(A[17]), .Q(n92) );
  NOR21 U453 ( .A(A[22]), .B(A[23]), .Q(n83) );
  NOR21 U454 ( .A(A[22]), .B(n95), .Q(n88) );
  NOR24 U455 ( .A(n398), .B(A[14]), .Q(n155) );
  NAND21 U456 ( .A(n110), .B(n96), .Q(n95) );
  INV1 U457 ( .A(n95), .Q(n93) );
  XNR21 U458 ( .A(A[22]), .B(n91), .Q(DIFF[22]) );
  OAI212 U459 ( .A(n195), .B(n191), .C(n192), .Q(n186) );
  OAI212 U460 ( .A(n176), .B(n372), .C(n177), .Q(n175) );
  OAI212 U461 ( .A(n202), .B(n210), .C(n203), .Q(n201) );
  NOR24 U462 ( .A(n401), .B(A[16]), .Q(n135) );
  NOR24 U463 ( .A(n395), .B(A[15]), .Q(n142) );
  CLKIN0 U464 ( .A(B[6]), .Q(n259) );
  OAI211 U465 ( .A(n393), .B(n391), .C(n88), .Q(n86) );
  XNR22 U466 ( .A(A[26]), .B(n63), .Q(DIFF[26]) );
  OAI212 U467 ( .A(n394), .B(n391), .C(n110), .Q(n104) );
  OAI212 U468 ( .A(n158), .B(n372), .C(n159), .Q(n157) );
  XNR22 U469 ( .A(A[27]), .B(n56), .Q(DIFF[27]) );
  OAI212 U470 ( .A(n166), .B(n131), .C(n132), .Q(n130) );
  NOR21 U471 ( .A(A[24]), .B(n79), .Q(n72) );
  NAND26 U472 ( .A(A[13]), .B(n397), .Q(n163) );
  AOI212 U473 ( .A(n197), .B(n129), .C(n130), .Q(n2) );
  NAND22 U474 ( .A(n238), .B(n163), .Q(n21) );
  CLKIN3 U475 ( .A(n163), .Q(n161) );
  NAND20 U476 ( .A(n244), .B(n210), .Q(n27) );
  NOR24 U477 ( .A(n379), .B(n223), .Q(n212) );
  INV3 U478 ( .A(B[4]), .Q(n404) );
  NAND22 U479 ( .A(n167), .B(n238), .Q(n158) );
  INV0 U480 ( .A(B[8]), .Q(n257) );
  XNR21 U481 ( .A(A[20]), .B(n104), .Q(DIFF[20]) );
  INV3 U482 ( .A(n108), .Q(n110) );
  CLKIN0 U483 ( .A(n67), .Q(n66) );
  NAND20 U484 ( .A(n241), .B(n192), .Q(n24) );
  XNR21 U485 ( .A(n29), .B(n225), .Q(DIFF[5]) );
  NOR21 U486 ( .A(n59), .B(n49), .Q(n48) );
  NOR20 U487 ( .A(n47), .B(n34), .Q(n33) );
  NAND20 U488 ( .A(n185), .B(n240), .Q(n176) );
  AOI212 U489 ( .A(n247), .B(n231), .C(n228), .Q(n226) );
  XNR20 U490 ( .A(A[3]), .B(A[2]), .Q(DIFF[3]) );
  INV0 U491 ( .A(A[2]), .Q(DIFF[2]) );
  NOR20 U492 ( .A(A[3]), .B(A[2]), .Q(n3) );
  INV3 U493 ( .A(n162), .Q(n238) );
  INV3 U494 ( .A(n59), .Q(n60) );
  INV3 U495 ( .A(B[7]), .Q(n403) );
  NAND22 U496 ( .A(n96), .B(n83), .Q(n82) );
  INV0 U497 ( .A(A[28]), .Q(n50) );
  AOI211 U498 ( .A(n168), .B(n140), .C(n141), .Q(n139) );
  INV3 U499 ( .A(n392), .Q(n394) );
  INV3 U500 ( .A(n35), .Q(n34) );
  NOR20 U501 ( .A(A[29]), .B(A[30]), .Q(n35) );
  INV3 U502 ( .A(B[5]), .Q(n405) );
  INV0 U503 ( .A(n135), .Q(n235) );
  INV0 U504 ( .A(n155), .Q(n237) );
  NOR20 U505 ( .A(A[18]), .B(n125), .Q(n118) );
  NOR20 U506 ( .A(A[20]), .B(n108), .Q(n101) );
  NOR21 U507 ( .A(n66), .B(n79), .Q(n65) );
  NOR20 U508 ( .A(A[29]), .B(n47), .Q(n40) );
  INV3 U509 ( .A(B[12]), .Q(n400) );
  INV3 U510 ( .A(B[13]), .Q(n397) );
  INV3 U511 ( .A(B[14]), .Q(n398) );
  INV3 U512 ( .A(B[16]), .Q(n401) );
  AOI211 U513 ( .A(n205), .B(n225), .C(n206), .Q(n204) );
  INV3 U514 ( .A(B[10]), .Q(n399) );
  INV3 U515 ( .A(B[11]), .Q(n254) );
  INV3 U516 ( .A(B[15]), .Q(n395) );
  INV3 U517 ( .A(B[17]), .Q(n402) );
  XOR21 U518 ( .A(n26), .B(n204), .Q(DIFF[8]) );
  XNR21 U519 ( .A(n231), .B(n30), .Q(DIFF[4]) );
  NAND22 U520 ( .A(n247), .B(n230), .Q(n30) );
  BUF2 U521 ( .A(A[0]), .Q(DIFF[0]) );
  BUF2 U522 ( .A(A[1]), .Q(DIFF[1]) );
  CLKIN3 U523 ( .A(n3), .Q(n231) );
  AOI211 U524 ( .A(n225), .B(n368), .C(n363), .Q(n211) );
endmodule


module sqroot_comb_NBITS32_DW01_inc_3 ( A, SUM );
  input [16:0] A;
  output [16:0] SUM;
  wire   n1, n2, n3, n6, n7, n9, n10, n11, n12, n14, n15, n17, n18, n19, n21,
         n24, n25, n26, n27, n29, n30, n31, n32, n33, n36, n37, n38, n39, n41,
         n42, n44, n45, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57,
         n58, n59, n60, n62, n63, n64, n69, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n128, n129, n130;

  CLKIN1 U97 ( .A(A[0]), .Q(SUM[0]) );
  CLKIN0 U98 ( .A(A[3]), .Q(n130) );
  NAND22 U99 ( .A(n63), .B(n57), .Q(n56) );
  NAND21 U100 ( .A(n63), .B(n47), .Q(n46) );
  NOR21 U101 ( .A(n130), .B(n64), .Q(n60) );
  NAND22 U102 ( .A(n7), .B(A[15]), .Q(n3) );
  INV2 U103 ( .A(n3), .Q(n2) );
  INV0 U104 ( .A(A[13]), .Q(n116) );
  INV1 U105 ( .A(n56), .Q(n55) );
  INV2 U106 ( .A(n1), .Q(SUM[16]) );
  INV6 U107 ( .A(SUM[0]), .Q(n125) );
  CLKIN1 U108 ( .A(SUM[0]), .Q(n126) );
  CLKIN0 U109 ( .A(A[1]), .Q(n128) );
  NOR20 U110 ( .A(n21), .B(n128), .Q(n18) );
  CLKIN0 U111 ( .A(A[2]), .Q(n129) );
  CLKIN0 U112 ( .A(n27), .Q(n26) );
  INV0 U113 ( .A(n48), .Q(n47) );
  INV0 U114 ( .A(A[10]), .Q(n121) );
  INV0 U115 ( .A(A[12]), .Q(n119) );
  CLKIN0 U116 ( .A(A[4]), .Q(n58) );
  NAND20 U117 ( .A(n125), .B(n63), .Q(n62) );
  NAND20 U118 ( .A(n125), .B(n60), .Q(n59) );
  XNR20 U119 ( .A(A[9]), .B(n36), .Q(SUM[9]) );
  NAND20 U120 ( .A(n125), .B(n52), .Q(n51) );
  NAND20 U121 ( .A(n125), .B(n55), .Q(n54) );
  NAND20 U122 ( .A(n125), .B(n30), .Q(n29) );
  NAND20 U123 ( .A(n125), .B(n18), .Q(n17) );
  INV3 U124 ( .A(A[7]), .Q(n117) );
  NOR21 U125 ( .A(n129), .B(n128), .Q(n63) );
  INV3 U126 ( .A(n63), .Q(n64) );
  INV3 U127 ( .A(n18), .Q(n19) );
  INV3 U128 ( .A(A[5]), .Q(n124) );
  NAND22 U129 ( .A(n27), .B(A[11]), .Q(n21) );
  NOR21 U130 ( .A(n122), .B(n11), .Q(n7) );
  NOR21 U131 ( .A(n38), .B(n46), .Q(n37) );
  INV3 U132 ( .A(n39), .Q(n38) );
  NOR20 U133 ( .A(n31), .B(n128), .Q(n30) );
  NAND22 U134 ( .A(n18), .B(n12), .Q(n11) );
  NOR21 U135 ( .A(n116), .B(n119), .Q(n12) );
  NOR21 U136 ( .A(n121), .B(n31), .Q(n27) );
  NOR21 U137 ( .A(n120), .B(n117), .Q(n39) );
  INV3 U138 ( .A(A[11]), .Q(n118) );
  INV3 U139 ( .A(A[14]), .Q(n122) );
  NOR21 U140 ( .A(n58), .B(n130), .Q(n57) );
  NAND20 U141 ( .A(A[2]), .B(n32), .Q(n31) );
  NOR21 U142 ( .A(n33), .B(n48), .Q(n32) );
  NAND22 U143 ( .A(n39), .B(A[9]), .Q(n33) );
  NAND22 U144 ( .A(n57), .B(n49), .Q(n48) );
  NOR21 U145 ( .A(n50), .B(n124), .Q(n49) );
  INV3 U146 ( .A(A[8]), .Q(n120) );
  INV3 U147 ( .A(A[15]), .Q(n123) );
  INV0 U148 ( .A(A[6]), .Q(n50) );
  XOR21 U149 ( .A(n121), .B(n29), .Q(SUM[10]) );
  XOR21 U150 ( .A(n123), .B(n6), .Q(SUM[15]) );
  NAND22 U151 ( .A(n126), .B(n7), .Q(n6) );
  XOR21 U152 ( .A(n58), .B(n59), .Q(SUM[4]) );
  XOR21 U153 ( .A(n130), .B(n62), .Q(SUM[3]) );
  XOR21 U154 ( .A(n119), .B(n17), .Q(SUM[12]) );
  XOR21 U155 ( .A(n129), .B(n69), .Q(SUM[2]) );
  NAND20 U156 ( .A(n125), .B(A[1]), .Q(n69) );
  NAND20 U157 ( .A(n125), .B(n2), .Q(n1) );
  XOR21 U158 ( .A(n124), .B(n54), .Q(SUM[5]) );
  XOR21 U159 ( .A(n116), .B(n14), .Q(SUM[13]) );
  NAND22 U160 ( .A(n125), .B(n15), .Q(n14) );
  NOR21 U161 ( .A(n119), .B(n19), .Q(n15) );
  XOR21 U162 ( .A(n117), .B(n44), .Q(SUM[7]) );
  NAND22 U163 ( .A(n125), .B(n45), .Q(n44) );
  INV3 U164 ( .A(n46), .Q(n45) );
  XOR21 U165 ( .A(n50), .B(n51), .Q(SUM[6]) );
  NOR21 U166 ( .A(n124), .B(n56), .Q(n52) );
  XOR21 U167 ( .A(n120), .B(n41), .Q(SUM[8]) );
  NAND22 U168 ( .A(n125), .B(n42), .Q(n41) );
  NOR21 U169 ( .A(n117), .B(n46), .Q(n42) );
  NAND22 U170 ( .A(n125), .B(n37), .Q(n36) );
  XOR21 U171 ( .A(n118), .B(n24), .Q(SUM[11]) );
  NAND22 U172 ( .A(n125), .B(n25), .Q(n24) );
  NOR20 U173 ( .A(n26), .B(n128), .Q(n25) );
  XOR21 U174 ( .A(n122), .B(n9), .Q(SUM[14]) );
  NAND22 U175 ( .A(n126), .B(n10), .Q(n9) );
  INV1 U176 ( .A(n11), .Q(n10) );
  XNR21 U177 ( .A(n128), .B(n126), .Q(SUM[1]) );
endmodule


module sqroot_comb_NBITS32_DW01_sub_31 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n39, n40, n41,
         n44, n45, n46, n47, n51, n52, n53, n56, n57, n58, n60, n63, n64, n65,
         n68, n69, n70, n75, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n91, n92, n93, n94, n95, n96, n99, n100, n102, n103, n104, n105, n106,
         n107, n108, n109, n111, n114, n115, n116, n117, n118, n124, n125,
         n126, n127, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n139, n141, n142, n143, n144, n148, n149, n150, n151, n152, n153,
         n155, n158, n159, n160, n161, n163, n164, n165, n166, n168, n169,
         n170, n171, n172, n177, n178, n179, n180, n181, n182, n184, n185,
         n186, n187, n194, n197, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319;

  XOR22 U3 ( .A(A[30]), .B(n29), .Q(DIFF[30]) );
  NOR24 U18 ( .A(n57), .B(n35), .Q(n34) );
  XOR22 U24 ( .A(A[27]), .B(n44), .Q(DIFF[27]) );
  OAI212 U78 ( .A(n79), .B(n133), .C(n80), .Q(n1) );
  XOR22 U87 ( .A(n13), .B(n92), .Q(DIFF[19]) );
  XOR22 U97 ( .A(n105), .B(n14), .Q(DIFF[18]) );
  OAI212 U104 ( .A(n99), .B(n294), .C(n100), .Q(n94) );
  AOI212 U106 ( .A(n179), .B(n111), .C(n102), .Q(n100) );
  XOR22 U113 ( .A(n15), .B(n114), .Q(DIFF[17]) );
  NOR24 U123 ( .A(n314), .B(A[17]), .Q(n108) );
  AOI212 U126 ( .A(n132), .B(n115), .C(n116), .Q(n114) );
  AOI212 U134 ( .A(n181), .B(n129), .C(n124), .Q(n118) );
  XNR22 U149 ( .A(n18), .B(n142), .Q(DIFF[14]) );
  AOI212 U151 ( .A(n159), .B(n134), .C(n135), .Q(n133) );
  OAI212 U153 ( .A(n153), .B(n136), .C(n137), .Q(n135) );
  AOI212 U155 ( .A(n296), .B(n148), .C(n139), .Q(n137) );
  XNR22 U162 ( .A(n19), .B(n151), .Q(DIFF[13]) );
  OAI212 U163 ( .A(n143), .B(n158), .C(n144), .Q(n142) );
  OAI212 U186 ( .A(n172), .B(n160), .C(n161), .Q(n159) );
  AOI212 U188 ( .A(n168), .B(n186), .C(n163), .Q(n161) );
  NOR24 U205 ( .A(A[9]), .B(A[8]), .Q(n172) );
  NOR22 U226 ( .A(A[25]), .B(A[26]), .Q(n46) );
  INV0 U227 ( .A(n168), .Q(n293) );
  NOR22 U228 ( .A(n311), .B(A[18]), .Q(n103) );
  INV10 U229 ( .A(A[14]), .Q(n297) );
  INV8 U230 ( .A(n133), .Q(n132) );
  INV12 U231 ( .A(n108), .Q(n180) );
  NOR23 U232 ( .A(A[21]), .B(n310), .Q(n75) );
  NAND24 U233 ( .A(n93), .B(n81), .Q(n79) );
  NAND22 U234 ( .A(A[12]), .B(n312), .Q(n153) );
  NAND26 U235 ( .A(n179), .B(n180), .Q(n99) );
  NAND23 U236 ( .A(A[14]), .B(n194), .Q(n141) );
  XOR22 U237 ( .A(n12), .B(n85), .Q(DIFF[20]) );
  NOR22 U238 ( .A(n317), .B(A[19]), .Q(n88) );
  NOR23 U239 ( .A(A[23]), .B(A[24]), .Q(n60) );
  INV3 U240 ( .A(n172), .Q(n171) );
  INV8 U241 ( .A(n149), .Q(n184) );
  NAND21 U242 ( .A(A[16]), .B(n313), .Q(n126) );
  CLKIN2 U243 ( .A(B[12]), .Q(n312) );
  NOR23 U244 ( .A(n312), .B(A[12]), .Q(n152) );
  NAND24 U245 ( .A(A[10]), .B(n319), .Q(n170) );
  NAND28 U246 ( .A(n296), .B(n184), .Q(n136) );
  NAND28 U247 ( .A(B[14]), .B(n297), .Q(n296) );
  NOR24 U248 ( .A(n152), .B(n136), .Q(n134) );
  AOI212 U249 ( .A(n132), .B(n182), .C(n129), .Q(n127) );
  INV3 U250 ( .A(n88), .Q(n178) );
  INV3 U251 ( .A(n27), .Q(n26) );
  BUF2 U252 ( .A(A[7]), .Q(DIFF[7]) );
  INV0 U253 ( .A(A[8]), .Q(DIFF[8]) );
  NOR22 U254 ( .A(n33), .B(n310), .Q(n32) );
  AOI212 U255 ( .A(n181), .B(n129), .C(n124), .Q(n294) );
  CLKIN0 U256 ( .A(n118), .Q(n116) );
  NAND20 U257 ( .A(n187), .B(n293), .Q(n22) );
  XOR21 U258 ( .A(n20), .B(n158), .Q(DIFF[12]) );
  INV2 U259 ( .A(n159), .Q(n158) );
  NOR23 U260 ( .A(n52), .B(n310), .Q(n51) );
  NOR24 U261 ( .A(n197), .B(A[11]), .Q(n164) );
  INV3 U262 ( .A(n94), .Q(n96) );
  NAND23 U263 ( .A(A[11]), .B(n197), .Q(n165) );
  XOR21 U264 ( .A(A[29]), .B(n32), .Q(DIFF[29]) );
  NOR24 U265 ( .A(A[21]), .B(A[22]), .Q(n70) );
  NAND21 U266 ( .A(n58), .B(n46), .Q(n45) );
  NAND23 U267 ( .A(n187), .B(n186), .Q(n160) );
  NOR22 U268 ( .A(n30), .B(n310), .Q(n29) );
  NOR22 U269 ( .A(n45), .B(n310), .Q(n44) );
  CLKIN0 U270 ( .A(n83), .Q(n177) );
  NAND23 U271 ( .A(A[15]), .B(n316), .Q(n131) );
  INV4 U272 ( .A(n130), .Q(n182) );
  INV2 U273 ( .A(n96), .Q(n295) );
  XOR21 U274 ( .A(n21), .B(n166), .Q(DIFF[11]) );
  OAI212 U275 ( .A(n152), .B(n158), .C(n153), .Q(n151) );
  NOR22 U276 ( .A(n40), .B(n310), .Q(n39) );
  INV6 U277 ( .A(n164), .Q(n186) );
  CLKIN0 U278 ( .A(A[26]), .Q(n298) );
  NOR24 U279 ( .A(n57), .B(n310), .Q(n56) );
  NOR24 U280 ( .A(n64), .B(n310), .Q(n63) );
  INV3 U281 ( .A(n152), .Q(n185) );
  NAND21 U282 ( .A(A[19]), .B(n317), .Q(n91) );
  NOR23 U283 ( .A(n69), .B(n310), .Q(n68) );
  OAI211 U284 ( .A(n91), .B(n83), .C(n84), .Q(n82) );
  NOR23 U285 ( .A(n88), .B(n83), .Q(n81) );
  NAND20 U286 ( .A(n186), .B(n165), .Q(n21) );
  NOR22 U287 ( .A(A[28]), .B(A[27]), .Q(n36) );
  XOR22 U288 ( .A(A[31]), .B(n24), .Q(DIFF[31]) );
  NOR22 U289 ( .A(n25), .B(n310), .Q(n24) );
  NAND22 U290 ( .A(n34), .B(n26), .Q(n25) );
  INV1 U291 ( .A(A[29]), .Q(n31) );
  NOR20 U292 ( .A(A[27]), .B(n47), .Q(n41) );
  INV4 U293 ( .A(n126), .Q(n124) );
  INV2 U294 ( .A(n165), .Q(n163) );
  NOR24 U295 ( .A(n315), .B(A[13]), .Q(n149) );
  CLKIN0 U296 ( .A(B[11]), .Q(n197) );
  INV6 U297 ( .A(n57), .Q(n58) );
  NOR21 U298 ( .A(n313), .B(A[16]), .Q(n125) );
  NAND24 U299 ( .A(n300), .B(n301), .Q(DIFF[26]) );
  AOI211 U300 ( .A(n132), .B(n93), .C(n295), .Q(n92) );
  INV6 U301 ( .A(n170), .Q(n168) );
  XNR21 U302 ( .A(A[21]), .B(n310), .Q(DIFF[21]) );
  CLKIN3 U303 ( .A(n70), .Q(n69) );
  NAND24 U304 ( .A(n60), .B(n70), .Q(n57) );
  AOI212 U305 ( .A(n132), .B(n106), .C(n107), .Q(n105) );
  XOR22 U306 ( .A(A[28]), .B(n39), .Q(DIFF[28]) );
  NAND22 U307 ( .A(A[20]), .B(n318), .Q(n84) );
  XOR22 U308 ( .A(A[23]), .B(n68), .Q(DIFF[23]) );
  NAND26 U309 ( .A(A[17]), .B(n314), .Q(n109) );
  INV2 U310 ( .A(n34), .Q(n33) );
  XOR22 U311 ( .A(A[24]), .B(n63), .Q(DIFF[24]) );
  XOR22 U312 ( .A(A[22]), .B(n75), .Q(DIFF[22]) );
  CLKIN3 U313 ( .A(n93), .Q(n95) );
  NOR24 U314 ( .A(n99), .B(n117), .Q(n93) );
  NAND24 U315 ( .A(A[13]), .B(n315), .Q(n150) );
  INV6 U316 ( .A(n131), .Q(n129) );
  XOR22 U317 ( .A(A[25]), .B(n56), .Q(DIFF[25]) );
  NAND22 U318 ( .A(A[26]), .B(n299), .Q(n300) );
  NAND21 U319 ( .A(n298), .B(n51), .Q(n301) );
  CLKIN2 U320 ( .A(n51), .Q(n299) );
  XNR21 U321 ( .A(n17), .B(n132), .Q(DIFF[15]) );
  NAND21 U322 ( .A(n34), .B(n31), .Q(n30) );
  NOR23 U323 ( .A(n319), .B(A[10]), .Q(n169) );
  INV1 U324 ( .A(B[10]), .Q(n319) );
  OAI212 U325 ( .A(n88), .B(n96), .C(n91), .Q(n87) );
  NOR21 U326 ( .A(n88), .B(n95), .Q(n86) );
  NOR22 U327 ( .A(n316), .B(A[15]), .Q(n130) );
  INV3 U328 ( .A(n46), .Q(n47) );
  AOI211 U329 ( .A(n132), .B(n86), .C(n87), .Q(n85) );
  AOI212 U330 ( .A(n94), .B(n81), .C(n82), .Q(n80) );
  NAND22 U331 ( .A(n41), .B(n58), .Q(n40) );
  NAND20 U332 ( .A(n70), .B(n65), .Q(n64) );
  XNR21 U333 ( .A(n171), .B(n22), .Q(DIFF[10]) );
  CLKIN3 U334 ( .A(A[30]), .Q(n28) );
  INV0 U335 ( .A(n117), .Q(n115) );
  NOR24 U336 ( .A(n318), .B(A[20]), .Q(n83) );
  INV1 U337 ( .A(B[19]), .Q(n317) );
  NAND20 U338 ( .A(n184), .B(n150), .Q(n19) );
  INV0 U339 ( .A(B[14]), .Q(n194) );
  INV0 U340 ( .A(n153), .Q(n155) );
  INV3 U341 ( .A(n109), .Q(n111) );
  INV3 U342 ( .A(n104), .Q(n102) );
  NOR20 U343 ( .A(n108), .B(n117), .Q(n106) );
  NAND22 U344 ( .A(n58), .B(n53), .Q(n52) );
  CLKIN0 U345 ( .A(A[25]), .Q(n53) );
  NAND22 U346 ( .A(A[18]), .B(n311), .Q(n104) );
  NAND20 U347 ( .A(n177), .B(n84), .Q(n12) );
  INV3 U348 ( .A(n150), .Q(n148) );
  NAND22 U349 ( .A(n36), .B(n46), .Q(n35) );
  NAND24 U350 ( .A(n181), .B(n182), .Q(n117) );
  INV3 U351 ( .A(B[15]), .Q(n316) );
  INV3 U352 ( .A(B[16]), .Q(n313) );
  INV3 U353 ( .A(B[17]), .Q(n314) );
  NAND20 U354 ( .A(n178), .B(n91), .Q(n13) );
  NAND22 U355 ( .A(n28), .B(n31), .Q(n27) );
  INV3 U356 ( .A(A[23]), .Q(n65) );
  INV3 U357 ( .A(B[13]), .Q(n315) );
  INV3 U358 ( .A(B[18]), .Q(n311) );
  INV3 U359 ( .A(B[20]), .Q(n318) );
  INV3 U360 ( .A(n141), .Q(n139) );
  AOI210 U361 ( .A(n184), .B(n155), .C(n148), .Q(n144) );
  NAND20 U362 ( .A(n185), .B(n184), .Q(n143) );
  NAND20 U363 ( .A(n179), .B(n104), .Q(n14) );
  NAND20 U364 ( .A(n182), .B(n131), .Q(n17) );
  NAND20 U365 ( .A(n180), .B(n109), .Q(n15) );
  NAND20 U366 ( .A(n185), .B(n153), .Q(n20) );
  NAND20 U367 ( .A(n181), .B(n126), .Q(n16) );
  AOI210 U368 ( .A(n171), .B(n187), .C(n168), .Q(n166) );
  NAND20 U369 ( .A(n296), .B(n141), .Q(n18) );
  BUF2 U370 ( .A(A[5]), .Q(DIFF[5]) );
  BUF2 U371 ( .A(A[0]), .Q(DIFF[0]) );
  BUF2 U372 ( .A(A[1]), .Q(DIFF[1]) );
  BUF2 U373 ( .A(A[2]), .Q(DIFF[2]) );
  BUF2 U374 ( .A(A[3]), .Q(DIFF[3]) );
  BUF2 U375 ( .A(A[4]), .Q(DIFF[4]) );
  BUF6 U376 ( .A(A[6]), .Q(DIFF[6]) );
  XOR22 U377 ( .A(n16), .B(n127), .Q(DIFF[16]) );
  OAI210 U378 ( .A(n108), .B(n118), .C(n109), .Q(n107) );
  XNR20 U379 ( .A(A[9]), .B(A[8]), .Q(DIFF[9]) );
  BUF15 U380 ( .A(n1), .Q(n310) );
  CLKIN6 U381 ( .A(n169), .Q(n187) );
  CLKIN6 U382 ( .A(n125), .Q(n181) );
  CLKIN6 U383 ( .A(n103), .Q(n179) );
endmodule


module sqroot_comb_NBITS32_DW01_sub_32 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n12, n13, n14, n15, n16, n18, n19, n20, n21, n22, n23, n24,
         n27, n28, n29, n30, n32, n34, n35, n36, n39, n41, n42, n45, n47, n48,
         n49, n53, n55, n56, n59, n61, n63, n67, n70, n71, n72, n74, n76, n77,
         n78, n79, n80, n81, n84, n85, n86, n87, n88, n89, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n108, n110, n111,
         n112, n113, n114, n115, n119, n120, n121, n122, n123, n124, n125,
         n126, n130, n131, n132, n134, n135, n137, n140, n146, n147, n148,
         n151, n153, n156, n157, n158, n159, n162, n165, n166, n167, n168,
         n169, n170, n171, n178, n181, net715484, net715516, net715620,
         net716252, net720562, net722922, net724321, net724323, net716232, n17,
         n133, net725924, n154, n145, n143, n142, n152, n150, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n314, n315, n316, n317, n318, n319,
         n320;

  XOR22 U1 ( .A(A[31]), .B(n22), .Q(DIFF[31]) );
  XNR22 U14 ( .A(A[28]), .B(n314), .Q(DIFF[28]) );
  OAI212 U20 ( .A(n290), .B(n294), .C(n34), .Q(n1) );
  XOR22 U28 ( .A(A[26]), .B(n45), .Q(DIFF[26]) );
  AOI212 U104 ( .A(n103), .B(n99), .C(n100), .Q(n98) );
  AOI212 U113 ( .A(net724321), .B(n105), .C(n106), .Q(n104) );
  NOR24 U114 ( .A(n123), .B(n285), .Q(n105) );
  OAI212 U115 ( .A(n285), .B(n124), .C(n108), .Q(n106) );
  XNR22 U124 ( .A(n16), .B(n122), .Q(DIFF[17]) );
  AOI212 U143 ( .A(n137), .B(n167), .C(n130), .Q(n124) );
  XNR22 U136 ( .A(n17), .B(n133), .Q(DIFF[16]) );
  AOI212 U164 ( .A(n169), .B(n150), .C(n145), .Q(n143) );
  INV6 U207 ( .A(n134), .Q(n274) );
  INV1 U208 ( .A(n134), .Q(n168) );
  INV6 U209 ( .A(n120), .Q(n275) );
  INV1 U210 ( .A(n120), .Q(n166) );
  OAI210 U211 ( .A(net720562), .B(n151), .C(n152), .Q(net724323) );
  XOR21 U212 ( .A(A[23]), .B(n70), .Q(DIFF[23]) );
  INV3 U213 ( .A(B[12]), .Q(n181) );
  NAND22 U214 ( .A(A[16]), .B(net715484), .Q(n132) );
  NAND23 U215 ( .A(A[30]), .B(n277), .Q(n278) );
  NAND22 U216 ( .A(n276), .B(n27), .Q(n279) );
  NAND28 U217 ( .A(n278), .B(n279), .Q(DIFF[30]) );
  INV0 U218 ( .A(A[30]), .Q(n276) );
  CLKIN6 U219 ( .A(n27), .Q(n277) );
  CLKIN12 U220 ( .A(n96), .Q(n94) );
  NOR23 U221 ( .A(n318), .B(A[18]), .Q(n111) );
  NAND21 U222 ( .A(n166), .B(n289), .Q(n16) );
  INV1 U223 ( .A(net716252), .Q(n280) );
  INV1 U224 ( .A(n137), .Q(net716252) );
  NAND23 U225 ( .A(A[27]), .B(n282), .Q(n283) );
  NOR23 U226 ( .A(A[25]), .B(A[24]), .Q(n48) );
  AOI212 U227 ( .A(n287), .B(n79), .C(n80), .Q(n78) );
  NAND28 U228 ( .A(n275), .B(n165), .Q(n285) );
  CLKIN3 U229 ( .A(n103), .Q(n294) );
  NAND24 U230 ( .A(n77), .B(n84), .Q(n76) );
  NOR23 U231 ( .A(n23), .B(n314), .Q(n22) );
  NAND21 U232 ( .A(n169), .B(n147), .Q(n19) );
  NAND24 U233 ( .A(A[12]), .B(n181), .Q(n158) );
  CLKIN8 U234 ( .A(n146), .Q(n169) );
  NAND28 U235 ( .A(A[15]), .B(n178), .Q(n135) );
  XOR22 U236 ( .A(n293), .B(n78), .Q(DIFF[22]) );
  OAI211 U237 ( .A(n81), .B(n292), .C(n74), .Q(n72) );
  INV3 U238 ( .A(n113), .Q(n301) );
  NAND23 U239 ( .A(n32), .B(n29), .Q(n28) );
  NAND22 U240 ( .A(n302), .B(n303), .Q(DIFF[18]) );
  INV6 U241 ( .A(n157), .Q(n171) );
  AOI212 U242 ( .A(n287), .B(n71), .C(n55), .Q(n53) );
  NAND24 U243 ( .A(n13), .B(n296), .Q(n297) );
  NAND22 U244 ( .A(n39), .B(n281), .Q(n284) );
  NAND24 U245 ( .A(n283), .B(n284), .Q(DIFF[27]) );
  INV0 U246 ( .A(A[27]), .Q(n281) );
  CLKIN3 U247 ( .A(n39), .Q(n282) );
  INV0 U248 ( .A(n156), .Q(net722922) );
  NAND26 U249 ( .A(n297), .B(n298), .Q(DIFF[20]) );
  INV6 U250 ( .A(n61), .Q(n63) );
  OAI212 U251 ( .A(n81), .B(n89), .C(n67), .Q(n61) );
  INV3 U252 ( .A(n98), .Q(n296) );
  INV6 U253 ( .A(net725924), .Q(n140) );
  AOI211 U254 ( .A(n168), .B(net725924), .C(n280), .Q(net716232) );
  NAND22 U255 ( .A(n94), .B(n97), .Q(n13) );
  NAND24 U256 ( .A(n162), .B(n86), .Q(n290) );
  XNR21 U257 ( .A(n159), .B(n21), .Q(DIFF[12]) );
  INV3 U258 ( .A(n290), .Q(n79) );
  CLKIN3 U259 ( .A(net724323), .Q(n148) );
  INV6 U260 ( .A(n152), .Q(n150) );
  NAND24 U261 ( .A(A[13]), .B(net715620), .Q(n152) );
  CLKIN0 U262 ( .A(B[13]), .Q(net715620) );
  NAND20 U263 ( .A(n170), .B(n152), .Q(n20) );
  OAI212 U264 ( .A(n142), .B(n154), .C(n143), .Q(net725924) );
  NAND24 U265 ( .A(n170), .B(n169), .Q(n142) );
  AOI212 U266 ( .A(n171), .B(n159), .C(n156), .Q(n154) );
  INV3 U267 ( .A(n147), .Q(n145) );
  NAND22 U268 ( .A(A[14]), .B(net715516), .Q(n147) );
  OAI212 U269 ( .A(n142), .B(n154), .C(n143), .Q(net724321) );
  NAND20 U270 ( .A(n167), .B(n132), .Q(n17) );
  CLKIN10 U271 ( .A(n131), .Q(n167) );
  INV3 U272 ( .A(net716232), .Q(n133) );
  INV12 U273 ( .A(n135), .Q(n137) );
  OAI212 U274 ( .A(n81), .B(n89), .C(n67), .Q(n286) );
  NOR23 U275 ( .A(n320), .B(A[21]), .Q(n81) );
  NAND22 U276 ( .A(n125), .B(n166), .Q(n114) );
  INV2 U277 ( .A(n294), .Q(n287) );
  NOR24 U278 ( .A(net715484), .B(A[16]), .Q(n131) );
  AOI211 U279 ( .A(n315), .B(n86), .C(n87), .Q(n85) );
  INV6 U280 ( .A(n104), .Q(n103) );
  NOR23 U281 ( .A(net715516), .B(A[14]), .Q(n146) );
  NAND26 U282 ( .A(A[19]), .B(n316), .Q(n102) );
  NOR24 U283 ( .A(n76), .B(A[23]), .Q(n67) );
  XNR22 U284 ( .A(A[11]), .B(A[10]), .Q(DIFF[11]) );
  NOR22 U285 ( .A(n286), .B(n35), .Q(n34) );
  NOR24 U286 ( .A(net715620), .B(A[13]), .Q(n151) );
  NOR24 U287 ( .A(n181), .B(A[12]), .Q(n157) );
  NAND22 U288 ( .A(A[18]), .B(n318), .Q(n112) );
  INV3 U289 ( .A(A[22]), .Q(n77) );
  NOR22 U290 ( .A(n316), .B(A[19]), .Q(n101) );
  INV6 U291 ( .A(n88), .Q(n86) );
  INV2 U292 ( .A(net720562), .Q(n153) );
  INV2 U293 ( .A(n125), .Q(n288) );
  INV1 U294 ( .A(n123), .Q(n125) );
  INV0 U295 ( .A(n119), .Q(n289) );
  AOI211 U296 ( .A(n171), .B(n159), .C(n156), .Q(net720562) );
  AOI211 U297 ( .A(n137), .B(n167), .C(n130), .Q(n299) );
  NAND28 U298 ( .A(n274), .B(n167), .Q(n123) );
  INV6 U299 ( .A(n121), .Q(n119) );
  INV2 U300 ( .A(n48), .Q(n49) );
  XOR22 U301 ( .A(A[29]), .B(n30), .Q(DIFF[29]) );
  XOR22 U302 ( .A(n12), .B(n85), .Q(DIFF[21]) );
  CLKIN0 U303 ( .A(B[15]), .Q(n178) );
  CLKIN0 U304 ( .A(n77), .Q(n293) );
  NAND26 U305 ( .A(n99), .B(n94), .Q(n88) );
  INV1 U306 ( .A(n126), .Q(n291) );
  INV3 U307 ( .A(n299), .Q(n126) );
  AOI212 U308 ( .A(n94), .B(n100), .C(n95), .Q(n292) );
  INV1 U309 ( .A(A[29]), .Q(n29) );
  CLKBU15 U310 ( .A(n103), .Q(n315) );
  INV6 U311 ( .A(n158), .Q(n156) );
  NAND21 U312 ( .A(n63), .B(n48), .Q(n47) );
  NAND23 U313 ( .A(n63), .B(n42), .Q(n41) );
  NAND21 U314 ( .A(n63), .B(n56), .Q(n55) );
  INV2 U315 ( .A(n292), .Q(n87) );
  NAND22 U316 ( .A(n36), .B(n48), .Q(n35) );
  INV6 U317 ( .A(n111), .Q(n165) );
  NAND24 U318 ( .A(A[20]), .B(n319), .Q(n97) );
  INV6 U319 ( .A(n102), .Q(n100) );
  NAND22 U320 ( .A(n162), .B(n84), .Q(n12) );
  INV6 U321 ( .A(n132), .Q(n130) );
  CLKIN4 U322 ( .A(n97), .Q(n95) );
  NAND22 U323 ( .A(n295), .B(n98), .Q(n298) );
  INV1 U324 ( .A(n13), .Q(n295) );
  XOR21 U325 ( .A(n18), .B(n140), .Q(DIFF[15]) );
  INV3 U326 ( .A(A[28]), .Q(n32) );
  NAND22 U327 ( .A(n99), .B(n102), .Q(n14) );
  NOR24 U328 ( .A(n178), .B(A[15]), .Q(n134) );
  NOR24 U329 ( .A(n28), .B(n314), .Q(n27) );
  NOR21 U330 ( .A(A[26]), .B(n49), .Q(n42) );
  NAND21 U331 ( .A(n15), .B(n113), .Q(n302) );
  AOI211 U332 ( .A(n166), .B(n126), .C(n119), .Q(n115) );
  NOR24 U333 ( .A(A[28]), .B(n314), .Q(n30) );
  XOR22 U334 ( .A(A[25]), .B(n53), .Q(DIFF[25]) );
  NOR24 U335 ( .A(n319), .B(A[20]), .Q(n96) );
  BUF15 U336 ( .A(n1), .Q(n314) );
  NAND24 U337 ( .A(n300), .B(n301), .Q(n303) );
  INV2 U338 ( .A(n15), .Q(n300) );
  NOR22 U339 ( .A(A[30]), .B(n28), .Q(n24) );
  AOI212 U340 ( .A(n119), .B(n165), .C(n110), .Q(n108) );
  NOR21 U341 ( .A(A[26]), .B(A[27]), .Q(n36) );
  OAI212 U342 ( .A(n114), .B(n140), .C(n115), .Q(n113) );
  AOI211 U343 ( .A(n103), .B(n71), .C(n286), .Q(n59) );
  NAND22 U344 ( .A(A[21]), .B(n320), .Q(n84) );
  XNR21 U345 ( .A(n14), .B(n103), .Q(DIFF[19]) );
  XOR22 U346 ( .A(A[24]), .B(n59), .Q(DIFF[24]) );
  NOR24 U347 ( .A(n81), .B(n88), .Q(n71) );
  AOI212 U348 ( .A(n315), .B(n71), .C(n41), .Q(n39) );
  AOI212 U349 ( .A(n94), .B(n100), .C(n95), .Q(n89) );
  AOI211 U350 ( .A(n315), .B(n71), .C(n47), .Q(n45) );
  NOR24 U351 ( .A(n317), .B(A[17]), .Q(n120) );
  NAND23 U352 ( .A(A[17]), .B(n317), .Q(n121) );
  INV0 U353 ( .A(A[24]), .Q(n56) );
  INV0 U354 ( .A(n76), .Q(n74) );
  INV2 U355 ( .A(n24), .Q(n23) );
  XNR20 U356 ( .A(n20), .B(n153), .Q(DIFF[13]) );
  INV3 U357 ( .A(n81), .Q(n162) );
  INV3 U358 ( .A(B[16]), .Q(net715484) );
  INV3 U359 ( .A(B[17]), .Q(n317) );
  INV3 U360 ( .A(B[18]), .Q(n318) );
  INV3 U361 ( .A(B[20]), .Q(n319) );
  INV3 U362 ( .A(n112), .Q(n110) );
  INV3 U363 ( .A(B[14]), .Q(net715516) );
  INV3 U364 ( .A(B[19]), .Q(n316) );
  INV3 U365 ( .A(B[21]), .Q(n320) );
  NAND20 U366 ( .A(n165), .B(n112), .Q(n15) );
  INV3 U367 ( .A(n101), .Q(n99) );
  NAND20 U368 ( .A(n168), .B(net716252), .Q(n18) );
  XOR21 U369 ( .A(n19), .B(n148), .Q(DIFF[14]) );
  NAND20 U370 ( .A(n171), .B(net722922), .Q(n21) );
  INV3 U371 ( .A(n2), .Q(n159) );
  NOR21 U372 ( .A(A[11]), .B(A[10]), .Q(n2) );
  INV3 U373 ( .A(A[10]), .Q(DIFF[10]) );
  BUF2 U374 ( .A(A[0]), .Q(DIFF[0]) );
  BUF2 U375 ( .A(A[1]), .Q(DIFF[1]) );
  BUF2 U376 ( .A(A[2]), .Q(DIFF[2]) );
  BUF2 U377 ( .A(A[3]), .Q(DIFF[3]) );
  BUF2 U378 ( .A(A[4]), .Q(DIFF[4]) );
  BUF2 U379 ( .A(A[5]), .Q(DIFF[5]) );
  BUF2 U380 ( .A(A[6]), .Q(DIFF[6]) );
  BUF2 U381 ( .A(A[7]), .Q(DIFF[7]) );
  BUF2 U382 ( .A(A[8]), .Q(DIFF[8]) );
  BUF2 U383 ( .A(A[9]), .Q(DIFF[9]) );
  OAI212 U384 ( .A(n140), .B(n288), .C(n291), .Q(n122) );
  AOI212 U385 ( .A(n315), .B(n71), .C(n72), .Q(n70) );
  OAI210 U386 ( .A(n81), .B(n89), .C(n84), .Q(n80) );
  CLKIN6 U387 ( .A(n151), .Q(n170) );
endmodule


module sqroot_comb_NBITS32_DW01_sub_39 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n26,
         n27, n28, n29, n30, n31, n32, n33, n36, n37, n40, n41, n42, n45, n46,
         n47, n49, n50, n51, n52, n53, n54, n57, n58, n59, n61, n62, n65, n67,
         n69, n70, n75, n76, n77, n79, n80, n83, n85, n87, n89, n92, n95, n97,
         n98, n99, n100, n103, n104, n105, n107, n109, n114, n115, n116, n117,
         n118, n121, n122, n123, n124, n125, n126, n127, n129, n130, n131,
         n132, n133, n134, n135, n136, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n160, n161, n162, n163, n164, n165, n168, n169, n170, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n194, n195, n196, n197, n198, n199, n201,
         n202, n203, n204, n211, n214, n216, n313, n314, n315, n316, n317,
         n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
         n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
         n340, n341, n342, n343, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359;

  AOI212 U123 ( .A(n136), .B(n121), .C(n122), .Q(n116) );
  OAI212 U125 ( .A(n131), .B(n123), .C(n124), .Q(n122) );
  OAI212 U131 ( .A(n146), .B(n126), .C(n127), .Q(n125) );
  OAI212 U141 ( .A(n321), .B(n133), .C(n134), .Q(n132) );
  OAI212 U149 ( .A(n145), .B(n141), .C(n142), .Q(n136) );
  OAI212 U155 ( .A(n144), .B(n146), .C(n145), .Q(n143) );
  OAI212 U162 ( .A(n176), .B(n148), .C(n149), .Q(n147) );
  AOI212 U164 ( .A(n163), .B(n150), .C(n151), .Q(n149) );
  OAI212 U166 ( .A(n160), .B(n152), .C(n153), .Q(n151) );
  NOR24 U169 ( .A(n356), .B(A[14]), .Q(n152) );
  OAI212 U188 ( .A(n174), .B(n168), .C(n169), .Q(n163) );
  NOR24 U191 ( .A(n355), .B(A[12]), .Q(n168) );
  AOI212 U203 ( .A(n185), .B(n177), .C(n178), .Q(n176) );
  OAI212 U205 ( .A(n183), .B(n327), .C(n180), .Q(n178) );
  OAI212 U218 ( .A(n186), .B(n188), .C(n187), .Q(n185) );
  NAND24 U246 ( .A(n337), .B(n336), .Q(n339) );
  BUF2 U247 ( .A(n174), .Q(n313) );
  CLKIN4 U248 ( .A(n125), .Q(n333) );
  NOR23 U249 ( .A(n352), .B(A[11]), .Q(n173) );
  NAND23 U250 ( .A(n117), .B(n98), .Q(n58) );
  NAND23 U251 ( .A(n117), .B(n98), .Q(n76) );
  CLKIN3 U252 ( .A(n143), .Q(n337) );
  NAND23 U253 ( .A(n143), .B(n16), .Q(n338) );
  OAI212 U254 ( .A(n115), .B(n146), .C(n116), .Q(n114) );
  NOR23 U255 ( .A(n354), .B(A[16]), .Q(n141) );
  AOI211 U256 ( .A(n118), .B(n98), .C(n79), .Q(n77) );
  INV8 U257 ( .A(n51), .Q(n98) );
  NAND22 U258 ( .A(n117), .B(n98), .Q(n104) );
  NAND24 U259 ( .A(n92), .B(n109), .Q(n87) );
  NOR21 U260 ( .A(n42), .B(n32), .Q(n31) );
  NOR23 U261 ( .A(n87), .B(n53), .Q(n52) );
  NAND22 U262 ( .A(n54), .B(n70), .Q(n53) );
  NOR23 U263 ( .A(n358), .B(A[19]), .Q(n51) );
  INV6 U264 ( .A(n342), .Q(n343) );
  CLKIN6 U265 ( .A(n168), .Q(n342) );
  INV2 U266 ( .A(n70), .Q(n350) );
  NAND24 U267 ( .A(A[13]), .B(n211), .Q(n160) );
  INV0 U268 ( .A(n186), .Q(n204) );
  AOI212 U269 ( .A(n175), .B(n155), .C(n156), .Q(n154) );
  NAND23 U270 ( .A(n341), .B(n37), .Q(n36) );
  BUF2 U271 ( .A(A[4]), .Q(DIFF[4]) );
  BUF2 U272 ( .A(A[5]), .Q(DIFF[5]) );
  XOR21 U273 ( .A(n161), .B(n19), .Q(DIFF[13]) );
  INV3 U274 ( .A(B[10]), .Q(n214) );
  NOR23 U275 ( .A(n214), .B(A[10]), .Q(n327) );
  NAND20 U276 ( .A(n100), .B(n109), .Q(n99) );
  INV0 U277 ( .A(n109), .Q(n107) );
  NAND26 U278 ( .A(n324), .B(n325), .Q(DIFF[17]) );
  INV3 U279 ( .A(n15), .Q(n323) );
  BUF2 U280 ( .A(A[3]), .Q(DIFF[3]) );
  INV2 U281 ( .A(n329), .Q(n184) );
  NOR22 U282 ( .A(n141), .B(n144), .Q(n135) );
  OAI210 U283 ( .A(n188), .B(n186), .C(n187), .Q(n329) );
  INV2 U284 ( .A(n165), .Q(n314) );
  INV1 U285 ( .A(n163), .Q(n165) );
  NAND24 U286 ( .A(A[11]), .B(n352), .Q(n174) );
  NAND21 U287 ( .A(A[18]), .B(n357), .Q(n124) );
  NOR24 U288 ( .A(n216), .B(A[8]), .Q(n186) );
  BUF2 U289 ( .A(A[7]), .Q(n315) );
  BUF2 U290 ( .A(A[6]), .Q(n316) );
  AOI211 U291 ( .A(n118), .B(n98), .C(n87), .Q(n85) );
  CLKIN6 U292 ( .A(n87), .Q(n89) );
  XNR22 U293 ( .A(A[21]), .B(n95), .Q(DIFF[21]) );
  NAND24 U294 ( .A(n20), .B(n318), .Q(n319) );
  NAND22 U295 ( .A(n170), .B(n317), .Q(n320) );
  NAND23 U296 ( .A(n319), .B(n320), .Q(DIFF[12]) );
  INV3 U297 ( .A(n20), .Q(n317) );
  INV4 U298 ( .A(n170), .Q(n318) );
  CLKIN0 U299 ( .A(n136), .Q(n134) );
  NAND28 U300 ( .A(n338), .B(n339), .Q(DIFF[16]) );
  INV2 U301 ( .A(n328), .Q(n321) );
  OAI211 U302 ( .A(n176), .B(n148), .C(n149), .Q(n328) );
  NOR23 U303 ( .A(n179), .B(n182), .Q(n177) );
  NAND23 U304 ( .A(n132), .B(n15), .Q(n324) );
  NAND26 U305 ( .A(n322), .B(n323), .Q(n325) );
  INV3 U306 ( .A(n132), .Q(n322) );
  NAND21 U307 ( .A(n195), .B(n131), .Q(n15) );
  INV1 U308 ( .A(A[27]), .Q(n45) );
  INV1 U309 ( .A(n157), .Q(n199) );
  INV8 U310 ( .A(n147), .Q(n146) );
  OAI211 U311 ( .A(n330), .B(n165), .C(n160), .Q(n156) );
  BUF2 U312 ( .A(n188), .Q(n326) );
  NOR24 U313 ( .A(n214), .B(A[10]), .Q(n179) );
  XOR21 U314 ( .A(A[26]), .B(n341), .Q(DIFF[26]) );
  XOR22 U315 ( .A(n100), .B(n103), .Q(DIFF[20]) );
  INV3 U316 ( .A(A[20]), .Q(n100) );
  OAI211 U317 ( .A(n104), .B(n146), .C(n105), .Q(n103) );
  NAND22 U318 ( .A(n341), .B(n27), .Q(n26) );
  NAND23 U319 ( .A(n341), .B(n41), .Q(n40) );
  NOR23 U320 ( .A(A[7]), .B(A[6]), .Q(n188) );
  XOR22 U321 ( .A(n18), .B(n154), .Q(DIFF[14]) );
  NOR21 U322 ( .A(n330), .B(n164), .Q(n155) );
  INV3 U323 ( .A(n199), .Q(n330) );
  NAND23 U324 ( .A(n341), .B(n47), .Q(n46) );
  XOR22 U325 ( .A(n331), .B(n114), .Q(DIFF[19]) );
  INV15 U326 ( .A(n13), .Q(n331) );
  NAND22 U327 ( .A(n342), .B(n169), .Q(n20) );
  INV2 U328 ( .A(n162), .Q(n164) );
  OAI212 U329 ( .A(n76), .B(n146), .C(n97), .Q(n95) );
  NOR24 U330 ( .A(n157), .B(n152), .Q(n150) );
  AOI211 U331 ( .A(n118), .B(n98), .C(n99), .Q(n97) );
  NAND26 U332 ( .A(n135), .B(n121), .Q(n115) );
  NAND22 U333 ( .A(A[8]), .B(n216), .Q(n187) );
  INV2 U334 ( .A(B[8]), .Q(n216) );
  NAND24 U335 ( .A(n162), .B(n150), .Q(n148) );
  NOR21 U336 ( .A(A[25]), .B(A[24]), .Q(n54) );
  NOR21 U337 ( .A(A[24]), .B(n350), .Q(n62) );
  NOR21 U338 ( .A(A[28]), .B(n42), .Q(n37) );
  NOR20 U339 ( .A(A[29]), .B(A[28]), .Q(n33) );
  OAI212 U340 ( .A(n51), .B(n116), .C(n52), .Q(n50) );
  XNR22 U341 ( .A(A[28]), .B(n40), .Q(DIFF[28]) );
  NOR24 U342 ( .A(n123), .B(n130), .Q(n121) );
  NAND24 U343 ( .A(A[9]), .B(n359), .Q(n183) );
  NOR21 U344 ( .A(A[21]), .B(A[20]), .Q(n92) );
  NAND22 U345 ( .A(n125), .B(n14), .Q(n334) );
  NAND24 U346 ( .A(n332), .B(n333), .Q(n335) );
  NAND24 U347 ( .A(n334), .B(n335), .Q(DIFF[18]) );
  INV3 U348 ( .A(n14), .Q(n332) );
  NAND21 U349 ( .A(n194), .B(n124), .Q(n14) );
  XNR22 U350 ( .A(A[22]), .B(n83), .Q(DIFF[22]) );
  XNR21 U351 ( .A(A[24]), .B(n65), .Q(DIFF[24]) );
  NAND21 U352 ( .A(n201), .B(n313), .Q(n21) );
  INV1 U353 ( .A(n16), .Q(n336) );
  NAND21 U354 ( .A(n196), .B(n142), .Q(n16) );
  INV0 U355 ( .A(n152), .Q(n198) );
  AOI212 U356 ( .A(n136), .B(n121), .C(n122), .Q(n340) );
  NAND21 U357 ( .A(A[16]), .B(n354), .Q(n142) );
  INV1 U358 ( .A(n141), .Q(n196) );
  INV2 U359 ( .A(n173), .Q(n201) );
  OAI211 U360 ( .A(n182), .B(n184), .C(n183), .Q(n181) );
  CLKIN0 U361 ( .A(n174), .Q(n172) );
  OAI211 U362 ( .A(n146), .B(n58), .C(n59), .Q(n57) );
  OAI211 U363 ( .A(n146), .B(n58), .C(n85), .Q(n83) );
  AOI212 U364 ( .A(n175), .B(n201), .C(n172), .Q(n170) );
  AOI210 U365 ( .A(n136), .B(n195), .C(n129), .Q(n127) );
  NAND21 U366 ( .A(A[14]), .B(n356), .Q(n153) );
  NAND22 U367 ( .A(n355), .B(A[12]), .Q(n169) );
  NAND20 U368 ( .A(n199), .B(n160), .Q(n19) );
  NOR24 U369 ( .A(n343), .B(n173), .Q(n162) );
  XNR21 U370 ( .A(A[31]), .B(n26), .Q(DIFF[31]) );
  NOR22 U371 ( .A(A[23]), .B(A[22]), .Q(n70) );
  XNR21 U372 ( .A(A[25]), .B(n57), .Q(DIFF[25]) );
  AOI211 U373 ( .A(n118), .B(n98), .C(n61), .Q(n59) );
  OAI211 U374 ( .A(n76), .B(n146), .C(n77), .Q(n75) );
  OAI211 U375 ( .A(n146), .B(n104), .C(n67), .Q(n65) );
  NAND21 U376 ( .A(n197), .B(n145), .Q(n17) );
  NAND26 U377 ( .A(A[15]), .B(n353), .Q(n145) );
  CLKBU15 U378 ( .A(n1), .Q(n341) );
  AOI212 U379 ( .A(n328), .B(n49), .C(n50), .Q(n1) );
  NAND26 U380 ( .A(A[17]), .B(n351), .Q(n131) );
  NOR24 U381 ( .A(n351), .B(A[17]), .Q(n130) );
  XNR22 U382 ( .A(A[29]), .B(n36), .Q(DIFF[29]) );
  NOR24 U383 ( .A(n353), .B(A[15]), .Q(n144) );
  XNR22 U384 ( .A(A[23]), .B(n75), .Q(DIFF[23]) );
  XNR22 U385 ( .A(A[27]), .B(n46), .Q(DIFF[27]) );
  INV6 U386 ( .A(n340), .Q(n118) );
  INV8 U387 ( .A(n115), .Q(n117) );
  AOI211 U388 ( .A(n118), .B(n98), .C(n69), .Q(n67) );
  NAND22 U389 ( .A(n98), .B(n109), .Q(n13) );
  NAND28 U390 ( .A(A[19]), .B(n358), .Q(n109) );
  NAND21 U391 ( .A(n341), .B(n31), .Q(n30) );
  AOI211 U392 ( .A(n175), .B(n162), .C(n314), .Q(n161) );
  NOR24 U393 ( .A(n211), .B(A[13]), .Q(n157) );
  NAND22 U394 ( .A(A[10]), .B(n214), .Q(n180) );
  NOR22 U395 ( .A(n51), .B(n115), .Q(n49) );
  INV3 U396 ( .A(n182), .Q(n203) );
  NOR24 U397 ( .A(n359), .B(A[9]), .Q(n182) );
  INV2 U398 ( .A(n176), .Q(n175) );
  INV0 U399 ( .A(B[12]), .Q(n355) );
  CLKIN0 U400 ( .A(A[30]), .Q(n29) );
  INV3 U401 ( .A(n28), .Q(n27) );
  NAND22 U402 ( .A(n89), .B(n70), .Q(n69) );
  XNR21 U403 ( .A(n22), .B(n181), .Q(DIFF[10]) );
  NAND20 U404 ( .A(n202), .B(n180), .Q(n22) );
  CLKIN0 U405 ( .A(B[11]), .Q(n352) );
  AOI211 U406 ( .A(n118), .B(n98), .C(n107), .Q(n105) );
  INV1 U407 ( .A(B[18]), .Q(n357) );
  NOR24 U408 ( .A(n357), .B(A[18]), .Q(n123) );
  CLKIN2 U409 ( .A(n33), .Q(n32) );
  INV0 U410 ( .A(B[13]), .Q(n211) );
  INV3 U411 ( .A(B[9]), .Q(n359) );
  INV3 U412 ( .A(n42), .Q(n41) );
  INV3 U413 ( .A(n135), .Q(n133) );
  INV3 U414 ( .A(n123), .Q(n194) );
  INV3 U415 ( .A(n131), .Q(n129) );
  INV3 U416 ( .A(n130), .Q(n195) );
  NAND22 U417 ( .A(n62), .B(n89), .Q(n61) );
  NAND22 U418 ( .A(n45), .B(n47), .Q(n42) );
  XNR21 U419 ( .A(A[30]), .B(n30), .Q(DIFF[30]) );
  INV3 U420 ( .A(A[26]), .Q(n47) );
  NAND21 U421 ( .A(n135), .B(n195), .Q(n126) );
  NAND22 U422 ( .A(n31), .B(n29), .Q(n28) );
  INV3 U423 ( .A(B[14]), .Q(n356) );
  INV3 U424 ( .A(B[15]), .Q(n353) );
  INV3 U425 ( .A(B[16]), .Q(n354) );
  XNR21 U426 ( .A(n21), .B(n175), .Q(DIFF[11]) );
  NAND22 U427 ( .A(n89), .B(n80), .Q(n79) );
  CLKIN0 U428 ( .A(A[22]), .Q(n80) );
  INV3 U429 ( .A(B[17]), .Q(n351) );
  INV3 U430 ( .A(B[19]), .Q(n358) );
  NAND20 U431 ( .A(n198), .B(n153), .Q(n18) );
  XOR21 U432 ( .A(n146), .B(n17), .Q(DIFF[15]) );
  INV0 U433 ( .A(n144), .Q(n197) );
  INV0 U434 ( .A(n179), .Q(n202) );
  XOR20 U435 ( .A(n326), .B(n24), .Q(DIFF[8]) );
  NAND20 U436 ( .A(n204), .B(n187), .Q(n24) );
  XOR21 U437 ( .A(n23), .B(n184), .Q(DIFF[9]) );
  NAND20 U438 ( .A(n203), .B(n183), .Q(n23) );
  CLKIN0 U439 ( .A(n316), .Q(DIFF[6]) );
  XNR20 U440 ( .A(n316), .B(n315), .Q(DIFF[7]) );
  BUF2 U441 ( .A(A[1]), .Q(DIFF[1]) );
  BUF2 U442 ( .A(A[0]), .Q(DIFF[0]) );
  BUF2 U443 ( .A(A[2]), .Q(DIFF[2]) );
endmodule


module sqroot_comb_NBITS32_DW01_sub_43 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n2, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45,
         n46, n47, n48, n51, n52, n55, n56, n57, n58, n61, n62, n65, n66, n67,
         n69, n70, n73, n74, n77, n78, n79, n80, n83, n84, n87, n89, n90, n92,
         n95, n96, n99, n100, n101, n105, n106, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n126, n127,
         n128, n129, n130, n131, n132, n133, n136, n137, n138, n139, n140,
         n142, n143, n144, n145, n146, n147, n148, n149, n152, n153, n154,
         n155, n156, n157, n158, n160, n161, n162, n163, n164, n165, n166,
         n167, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n191, n192, n193, n194,
         n195, n196, n199, n200, n201, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n243, n246, n248, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378;

  AOI212 U109 ( .A(n178), .B(n110), .C(n111), .Q(n2) );
  OAI212 U111 ( .A(n147), .B(n112), .C(n113), .Q(n111) );
  OAI212 U133 ( .A(n128), .B(n177), .C(n129), .Q(n127) );
  OAI212 U141 ( .A(n136), .B(n144), .C(n137), .Q(n131) );
  OAI212 U157 ( .A(n146), .B(n177), .C(n356), .Q(n145) );
  AOI212 U163 ( .A(n167), .B(n152), .C(n153), .Q(n147) );
  OAI212 U165 ( .A(n162), .B(n154), .C(n155), .Q(n153) );
  OAI212 U181 ( .A(n164), .B(n177), .C(n165), .Q(n163) );
  OAI212 U189 ( .A(n176), .B(n172), .C(n173), .Q(n167) );
  OAI212 U195 ( .A(n175), .B(n177), .C(n176), .Q(n174) );
  AOI212 U204 ( .A(n194), .B(n181), .C(n182), .Q(n180) );
  OAI212 U206 ( .A(n191), .B(n183), .C(n184), .Q(n182) );
  OAI212 U228 ( .A(n199), .B(n205), .C(n200), .Q(n194) );
  AOI212 U243 ( .A(n208), .B(n216), .C(n209), .Q(n207) );
  OAI212 U245 ( .A(n214), .B(n210), .C(n211), .Q(n209) );
  OAI212 U251 ( .A(n213), .B(n215), .C(n357), .Q(n212) );
  OAI212 U258 ( .A(n217), .B(n219), .C(n218), .Q(n216) );
  NAND23 U287 ( .A(n130), .B(n114), .Q(n112) );
  NAND23 U288 ( .A(A[2]), .B(n376), .Q(n218) );
  NAND21 U289 ( .A(A[10]), .B(n243), .Q(n173) );
  NAND22 U290 ( .A(A[5]), .B(n248), .Q(n205) );
  NAND22 U291 ( .A(n148), .B(n225), .Q(n139) );
  CLKIN6 U292 ( .A(n147), .Q(n149) );
  INV1 U293 ( .A(n100), .Q(n101) );
  NOR24 U294 ( .A(A[18]), .B(A[17]), .Q(n100) );
  CLKIN3 U295 ( .A(n166), .Q(n164) );
  NAND26 U296 ( .A(n152), .B(n166), .Q(n146) );
  NAND23 U297 ( .A(A[9]), .B(n371), .Q(n176) );
  XNR22 U298 ( .A(n17), .B(n118), .Q(DIFF[16]) );
  INV4 U299 ( .A(n146), .Q(n148) );
  BUF2 U300 ( .A(n191), .Q(n354) );
  NAND20 U301 ( .A(n227), .B(n162), .Q(n22) );
  INV2 U302 ( .A(B[8]), .Q(n368) );
  NAND23 U303 ( .A(n70), .B(n80), .Q(n69) );
  CLKIN3 U304 ( .A(n66), .Q(n67) );
  NAND22 U305 ( .A(n366), .B(n34), .Q(n33) );
  NAND22 U306 ( .A(A[6]), .B(n375), .Q(n200) );
  NAND23 U307 ( .A(n366), .B(n106), .Q(n105) );
  INV3 U308 ( .A(n23), .Q(n363) );
  INV0 U309 ( .A(n162), .Q(n160) );
  BUF2 U310 ( .A(n21), .Q(n355) );
  NAND22 U311 ( .A(n366), .B(n62), .Q(n61) );
  NAND22 U312 ( .A(n366), .B(n52), .Q(n51) );
  NOR23 U313 ( .A(n210), .B(n213), .Q(n208) );
  INV2 U314 ( .A(B[2]), .Q(n376) );
  INV6 U315 ( .A(n364), .Q(n365) );
  NAND24 U316 ( .A(n58), .B(n48), .Q(n47) );
  NOR22 U317 ( .A(A[28]), .B(A[27]), .Q(n48) );
  NAND26 U318 ( .A(n92), .B(n100), .Q(n89) );
  NOR24 U319 ( .A(n375), .B(A[6]), .Q(n199) );
  INV3 U320 ( .A(n358), .Q(n215) );
  NOR23 U321 ( .A(n372), .B(A[11]), .Q(n161) );
  OAI211 U322 ( .A(n139), .B(n177), .C(n140), .Q(n138) );
  AOI211 U323 ( .A(n149), .B(n225), .C(n142), .Q(n140) );
  NAND23 U324 ( .A(A[11]), .B(n372), .Q(n162) );
  NOR23 U325 ( .A(n188), .B(n183), .Q(n181) );
  AOI210 U326 ( .A(n121), .B(n149), .C(n122), .Q(n120) );
  OAI211 U327 ( .A(n123), .B(n133), .C(n126), .Q(n122) );
  NAND20 U328 ( .A(n214), .B(n235), .Q(n30) );
  NAND26 U329 ( .A(A[3]), .B(n377), .Q(n214) );
  INV2 U330 ( .A(n149), .Q(n356) );
  NAND26 U331 ( .A(n360), .B(n361), .Q(n362) );
  BUF2 U332 ( .A(n214), .Q(n357) );
  OAI211 U333 ( .A(n217), .B(n219), .C(n218), .Q(n358) );
  NAND21 U334 ( .A(A[16]), .B(n374), .Q(n117) );
  NAND21 U335 ( .A(n222), .B(n117), .Q(n17) );
  CLKIN1 U336 ( .A(n116), .Q(n222) );
  NOR23 U337 ( .A(n116), .B(n123), .Q(n114) );
  INV2 U338 ( .A(n231), .Q(n359) );
  INV1 U339 ( .A(n188), .Q(n231) );
  NOR23 U340 ( .A(n246), .B(A[7]), .Q(n188) );
  AOI212 U341 ( .A(n131), .B(n114), .C(n115), .Q(n113) );
  CLKIN3 U342 ( .A(n172), .Q(n228) );
  INV0 U343 ( .A(n167), .Q(n165) );
  NOR23 U344 ( .A(n175), .B(n172), .Q(n166) );
  XNR22 U345 ( .A(n18), .B(n127), .Q(DIFF[15]) );
  XNR22 U346 ( .A(n29), .B(n212), .Q(DIFF[4]) );
  INV2 U347 ( .A(n57), .Q(n56) );
  OAI212 U348 ( .A(n126), .B(n116), .C(n117), .Q(n115) );
  XNR22 U349 ( .A(A[26]), .B(n61), .Q(DIFF[26]) );
  NAND24 U350 ( .A(A[4]), .B(n378), .Q(n211) );
  NOR21 U351 ( .A(A[19]), .B(n101), .Q(n96) );
  XNR22 U352 ( .A(A[27]), .B(n55), .Q(DIFF[27]) );
  NOR22 U353 ( .A(A[27]), .B(n57), .Q(n52) );
  XNR21 U354 ( .A(A[28]), .B(n51), .Q(DIFF[28]) );
  NAND22 U355 ( .A(n366), .B(n74), .Q(n73) );
  NAND23 U356 ( .A(A[7]), .B(n246), .Q(n191) );
  BUF15 U357 ( .A(n2), .Q(n366) );
  INV6 U358 ( .A(n179), .Q(n361) );
  NAND24 U359 ( .A(n193), .B(n181), .Q(n179) );
  CLKIN6 U360 ( .A(n207), .Q(n360) );
  XNR22 U361 ( .A(A[19]), .B(n99), .Q(DIFF[19]) );
  NAND23 U362 ( .A(A[15]), .B(n373), .Q(n126) );
  CLKIN3 U363 ( .A(n136), .Q(n224) );
  NOR23 U364 ( .A(n143), .B(n136), .Q(n130) );
  XNR22 U365 ( .A(A[31]), .B(n33), .Q(DIFF[31]) );
  NAND21 U366 ( .A(n225), .B(n144), .Q(n20) );
  INV0 U367 ( .A(n144), .Q(n142) );
  NAND28 U368 ( .A(n362), .B(n180), .Q(n178) );
  INV15 U369 ( .A(n178), .Q(n177) );
  NAND22 U370 ( .A(n66), .B(n46), .Q(n45) );
  XOR22 U371 ( .A(n363), .B(n174), .Q(DIFF[10]) );
  CLKIN3 U372 ( .A(n123), .Q(n223) );
  NOR21 U373 ( .A(n123), .B(n132), .Q(n121) );
  NAND22 U374 ( .A(n366), .B(n40), .Q(n39) );
  NOR23 U375 ( .A(n146), .B(n112), .Q(n110) );
  OAI211 U376 ( .A(n177), .B(n119), .C(n120), .Q(n118) );
  NAND21 U377 ( .A(A[12]), .B(n369), .Q(n155) );
  NAND22 U378 ( .A(n366), .B(n66), .Q(n65) );
  NOR22 U379 ( .A(n199), .B(n204), .Q(n193) );
  INV0 U380 ( .A(n194), .Q(n196) );
  NAND22 U381 ( .A(n232), .B(n200), .Q(n27) );
  XOR21 U382 ( .A(n26), .B(n192), .Q(DIFF[7]) );
  NOR23 U383 ( .A(n154), .B(n161), .Q(n152) );
  XNR22 U384 ( .A(A[25]), .B(n65), .Q(DIFF[25]) );
  CLKIN2 U385 ( .A(n130), .Q(n132) );
  NAND22 U386 ( .A(n366), .B(n96), .Q(n95) );
  XNR22 U387 ( .A(n20), .B(n145), .Q(DIFF[13]) );
  NAND23 U388 ( .A(n366), .B(n78), .Q(n77) );
  XNR22 U389 ( .A(A[29]), .B(n43), .Q(DIFF[29]) );
  NOR24 U390 ( .A(n374), .B(A[16]), .Q(n116) );
  NOR24 U391 ( .A(n243), .B(A[10]), .Q(n172) );
  AOI212 U392 ( .A(n365), .B(n186), .C(n187), .Q(n185) );
  OAI211 U393 ( .A(n359), .B(n196), .C(n354), .Q(n187) );
  NOR24 U394 ( .A(n377), .B(A[3]), .Q(n213) );
  XOR22 U395 ( .A(n25), .B(n185), .Q(DIFF[8]) );
  XOR21 U396 ( .A(A[17]), .B(n366), .Q(DIFF[17]) );
  XNR21 U397 ( .A(n28), .B(n365), .Q(DIFF[5]) );
  NAND22 U398 ( .A(n66), .B(n36), .Q(n35) );
  XNR21 U399 ( .A(A[23]), .B(n77), .Q(DIFF[23]) );
  NAND24 U400 ( .A(n66), .B(n58), .Q(n57) );
  OAI212 U401 ( .A(n157), .B(n177), .C(n158), .Q(n156) );
  NOR24 U402 ( .A(n373), .B(A[15]), .Q(n123) );
  NAND20 U403 ( .A(n121), .B(n148), .Q(n119) );
  NAND22 U404 ( .A(A[14]), .B(n367), .Q(n137) );
  NOR24 U405 ( .A(A[1]), .B(A[0]), .Q(n219) );
  NOR22 U406 ( .A(n248), .B(A[5]), .Q(n204) );
  NAND22 U407 ( .A(n366), .B(n44), .Q(n43) );
  NAND22 U408 ( .A(n366), .B(n90), .Q(n87) );
  NOR22 U409 ( .A(A[25]), .B(n67), .Q(n62) );
  NOR24 U410 ( .A(A[22]), .B(A[21]), .Q(n80) );
  NOR24 U411 ( .A(n376), .B(A[2]), .Q(n217) );
  NOR21 U412 ( .A(A[21]), .B(n89), .Q(n84) );
  NOR24 U413 ( .A(n367), .B(A[14]), .Q(n136) );
  NAND22 U414 ( .A(A[13]), .B(n370), .Q(n144) );
  XNR22 U415 ( .A(n163), .B(n22), .Q(DIFF[11]) );
  XOR22 U416 ( .A(n27), .B(n201), .Q(DIFF[6]) );
  NAND22 U417 ( .A(n236), .B(n218), .Q(n31) );
  NOR24 U418 ( .A(n378), .B(A[4]), .Q(n210) );
  NAND23 U419 ( .A(n90), .B(n80), .Q(n79) );
  INV4 U420 ( .A(n89), .Q(n90) );
  XNR21 U421 ( .A(A[22]), .B(n83), .Q(DIFF[22]) );
  NAND22 U422 ( .A(n366), .B(n84), .Q(n83) );
  NOR24 U423 ( .A(n371), .B(A[9]), .Q(n175) );
  NOR22 U424 ( .A(A[26]), .B(A[25]), .Q(n58) );
  XNR22 U425 ( .A(n355), .B(n156), .Q(DIFF[12]) );
  NOR24 U426 ( .A(n89), .B(n69), .Q(n66) );
  AOI212 U427 ( .A(n365), .B(n233), .C(n203), .Q(n201) );
  INV2 U428 ( .A(n131), .Q(n133) );
  NOR24 U429 ( .A(n368), .B(A[8]), .Q(n183) );
  CLKIN0 U430 ( .A(n183), .Q(n230) );
  NAND22 U431 ( .A(n366), .B(n100), .Q(n99) );
  NAND22 U432 ( .A(n366), .B(n56), .Q(n55) );
  XOR20 U433 ( .A(n219), .B(n31), .Q(DIFF[2]) );
  AOI211 U434 ( .A(n365), .B(n193), .C(n194), .Q(n192) );
  CLKIN4 U435 ( .A(n360), .Q(n364) );
  NOR24 U436 ( .A(n369), .B(A[12]), .Q(n154) );
  NAND21 U437 ( .A(n233), .B(n205), .Q(n28) );
  INV6 U438 ( .A(n161), .Q(n227) );
  NOR22 U439 ( .A(n370), .B(A[13]), .Q(n143) );
  XNR21 U440 ( .A(A[21]), .B(n87), .Q(DIFF[21]) );
  XNR21 U441 ( .A(A[18]), .B(n105), .Q(DIFF[18]) );
  INV0 U442 ( .A(B[14]), .Q(n367) );
  XNR21 U443 ( .A(A[24]), .B(n73), .Q(DIFF[24]) );
  INV3 U444 ( .A(A[30]), .Q(n38) );
  INV3 U445 ( .A(A[29]), .Q(n42) );
  NAND20 U446 ( .A(n226), .B(n155), .Q(n21) );
  INV0 U447 ( .A(n154), .Q(n226) );
  INV2 U448 ( .A(n35), .Q(n34) );
  INV0 U449 ( .A(A[17]), .Q(n106) );
  NAND20 U450 ( .A(n166), .B(n227), .Q(n157) );
  NAND20 U451 ( .A(n229), .B(n176), .Q(n24) );
  CLKIN0 U452 ( .A(B[3]), .Q(n377) );
  INV0 U453 ( .A(B[13]), .Q(n370) );
  NOR20 U454 ( .A(n359), .B(n195), .Q(n186) );
  NAND20 U455 ( .A(n231), .B(n354), .Q(n26) );
  INV0 U456 ( .A(n204), .Q(n233) );
  INV0 U457 ( .A(n213), .Q(n235) );
  XNR20 U458 ( .A(A[0]), .B(A[1]), .Q(DIFF[1]) );
  XNR21 U459 ( .A(n19), .B(n138), .Q(DIFF[14]) );
  NOR21 U460 ( .A(A[24]), .B(A[23]), .Q(n70) );
  XNR21 U461 ( .A(A[20]), .B(n95), .Q(DIFF[20]) );
  INV3 U462 ( .A(n143), .Q(n225) );
  NOR21 U463 ( .A(A[20]), .B(A[19]), .Q(n92) );
  NOR21 U464 ( .A(n37), .B(n47), .Q(n36) );
  NAND22 U465 ( .A(n42), .B(n38), .Q(n37) );
  XNR21 U466 ( .A(A[30]), .B(n39), .Q(DIFF[30]) );
  NOR21 U467 ( .A(A[29]), .B(n45), .Q(n40) );
  INV3 U468 ( .A(n47), .Q(n46) );
  NOR21 U469 ( .A(A[23]), .B(n79), .Q(n74) );
  NAND22 U470 ( .A(n223), .B(n126), .Q(n18) );
  INV2 U471 ( .A(n79), .Q(n78) );
  INV3 U472 ( .A(n45), .Q(n44) );
  INV3 U473 ( .A(B[6]), .Q(n375) );
  AOI210 U474 ( .A(n167), .B(n227), .C(n160), .Q(n158) );
  NAND22 U475 ( .A(n148), .B(n130), .Q(n128) );
  AOI211 U476 ( .A(n149), .B(n130), .C(n131), .Q(n129) );
  INV3 U477 ( .A(n175), .Q(n229) );
  NAND22 U478 ( .A(n224), .B(n137), .Q(n19) );
  NAND22 U479 ( .A(n228), .B(n173), .Q(n23) );
  INV3 U480 ( .A(B[4]), .Q(n378) );
  XOR20 U481 ( .A(n177), .B(n24), .Q(DIFF[9]) );
  INV0 U482 ( .A(n199), .Q(n232) );
  NAND22 U483 ( .A(n234), .B(n211), .Q(n29) );
  INV3 U484 ( .A(n210), .Q(n234) );
  INV3 U485 ( .A(B[11]), .Q(n372) );
  INV3 U486 ( .A(B[12]), .Q(n369) );
  INV3 U487 ( .A(B[15]), .Q(n373) );
  NAND22 U488 ( .A(n230), .B(n184), .Q(n25) );
  INV3 U489 ( .A(n205), .Q(n203) );
  NAND22 U490 ( .A(A[8]), .B(n368), .Q(n184) );
  CLKIN0 U491 ( .A(n193), .Q(n195) );
  INV3 U492 ( .A(B[9]), .Q(n371) );
  INV3 U493 ( .A(B[10]), .Q(n243) );
  INV3 U494 ( .A(B[16]), .Q(n374) );
  CLKIN0 U495 ( .A(n217), .Q(n236) );
  CLKIN0 U496 ( .A(B[5]), .Q(n248) );
  INV0 U497 ( .A(B[7]), .Q(n246) );
  XOR20 U498 ( .A(n30), .B(n215), .Q(DIFF[3]) );
endmodule


module sqroot_comb_NBITS32_DW_cmp_45 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n27, n42, n66, net715654, net715586, n9, n8, n7, n63, n61, n60, n6,
         n59, n58, n57, n56, n55, n54, n53, n52, n51, n50, n5, n49, n48, n47,
         n46, n45, n44, n43, n41, n40, n4, n39, n38, n37, n36, n35, n33, n31,
         n29, n23, n21, n20, n19, n18, n17, n16, n15, n14, n13, n12, n11, n10,
         n1, n34, n32, n30, n28, n26, n25, n24, n22, n141, n142, n143, n144,
         n145, n146, n147, n148, n149;

  NOR24 U5 ( .A(n7), .B(n5), .Q(n4) );
  OAI212 U40 ( .A(n40), .B(n43), .C(n41), .Q(n39) );
  OAI212 U53 ( .A(n53), .B(n56), .C(n54), .Q(n52) );
  OAI212 U58 ( .A(n60), .B(n58), .C(n59), .Q(n57) );
  AOI212 U51 ( .A(n57), .B(n51), .C(n52), .Q(n50) );
  OAI212 U36 ( .A(n36), .B(n50), .C(n37), .Q(n35) );
  AOI212 U11 ( .A(n35), .B(n11), .C(n12), .Q(n10) );
  OAI212 U13 ( .A(n19), .B(n22), .C(n13), .Q(n12) );
  NOR24 U26 ( .A(n141), .B(B[18]), .Q(n25) );
  OAI212 U31 ( .A(n31), .B(n34), .C(n32), .Q(n30) );
  AOI212 U23 ( .A(n23), .B(n30), .C(n24), .Q(n22) );
  NOR24 U78 ( .A(n19), .B(n21), .Q(n11) );
  NAND22 U79 ( .A(B[11]), .B(n147), .Q(n49) );
  OAI211 U80 ( .A(n46), .B(n49), .C(n47), .Q(n45) );
  INV4 U81 ( .A(B[27]), .Q(n8) );
  NOR23 U82 ( .A(n25), .B(n27), .Q(n23) );
  NAND22 U83 ( .A(B[17]), .B(net715654), .Q(n28) );
  NOR23 U84 ( .A(n17), .B(n14), .Q(n13) );
  NOR21 U85 ( .A(n46), .B(n48), .Q(n44) );
  NAND26 U86 ( .A(n10), .B(n1), .Q(GE_LT_GT_LE) );
  NOR24 U87 ( .A(n142), .B(B[16]), .Q(n31) );
  NAND22 U88 ( .A(B[15]), .B(net715586), .Q(n34) );
  INV3 U89 ( .A(A[15]), .Q(net715586) );
  NAND21 U90 ( .A(B[16]), .B(n142), .Q(n32) );
  INV0 U91 ( .A(A[16]), .Q(n142) );
  OAI212 U92 ( .A(n28), .B(n25), .C(n26), .Q(n24) );
  INV2 U93 ( .A(A[17]), .Q(net715654) );
  NAND21 U94 ( .A(B[18]), .B(n141), .Q(n26) );
  INV3 U95 ( .A(A[18]), .Q(n141) );
  NAND22 U96 ( .A(n44), .B(n38), .Q(n36) );
  NOR22 U97 ( .A(n146), .B(B[12]), .Q(n46) );
  NOR21 U98 ( .A(n147), .B(B[11]), .Q(n48) );
  CLKIN3 U99 ( .A(A[11]), .Q(n147) );
  NOR23 U100 ( .A(n42), .B(n40), .Q(n38) );
  NOR21 U101 ( .A(B[7]), .B(B[6]), .Q(n60) );
  NOR22 U102 ( .A(n61), .B(B[8]), .Q(n58) );
  INV2 U103 ( .A(A[8]), .Q(n61) );
  NAND20 U104 ( .A(B[8]), .B(n61), .Q(n59) );
  NOR22 U105 ( .A(n53), .B(n55), .Q(n51) );
  NOR24 U106 ( .A(n63), .B(B[10]), .Q(n53) );
  NOR21 U107 ( .A(n143), .B(B[9]), .Q(n55) );
  INV3 U108 ( .A(A[9]), .Q(n143) );
  NAND21 U109 ( .A(B[9]), .B(n143), .Q(n56) );
  NAND21 U110 ( .A(B[10]), .B(n63), .Q(n54) );
  CLKIN0 U111 ( .A(A[10]), .Q(n63) );
  AOI212 U112 ( .A(n38), .B(n45), .C(n39), .Q(n37) );
  NAND20 U113 ( .A(B[12]), .B(n146), .Q(n47) );
  INV3 U114 ( .A(A[12]), .Q(n146) );
  NOR23 U115 ( .A(n145), .B(B[14]), .Q(n40) );
  NAND22 U116 ( .A(B[13]), .B(n66), .Q(n43) );
  INV0 U117 ( .A(A[13]), .Q(n66) );
  NAND21 U118 ( .A(B[14]), .B(n145), .Q(n41) );
  INV3 U119 ( .A(A[14]), .Q(n145) );
  NOR24 U120 ( .A(n144), .B(B[19]), .Q(n19) );
  NAND23 U121 ( .A(n23), .B(n29), .Q(n21) );
  NOR22 U122 ( .A(n33), .B(n31), .Q(n29) );
  NOR23 U123 ( .A(net715586), .B(B[15]), .Q(n33) );
  NAND24 U124 ( .A(n18), .B(n20), .Q(n17) );
  NOR23 U125 ( .A(B[20]), .B(B[21]), .Q(n18) );
  NAND23 U126 ( .A(B[19]), .B(n144), .Q(n20) );
  INV3 U127 ( .A(A[19]), .Q(n144) );
  NAND26 U128 ( .A(n15), .B(n16), .Q(n14) );
  NOR24 U129 ( .A(B[25]), .B(B[24]), .Q(n15) );
  NOR24 U130 ( .A(B[23]), .B(B[22]), .Q(n16) );
  INV6 U131 ( .A(n148), .Q(n1) );
  NAND26 U132 ( .A(n4), .B(n149), .Q(n148) );
  NAND24 U133 ( .A(n8), .B(n9), .Q(n7) );
  INV6 U134 ( .A(B[26]), .Q(n9) );
  INV6 U135 ( .A(n6), .Q(n5) );
  NOR24 U136 ( .A(B[29]), .B(B[28]), .Q(n6) );
  NOR24 U137 ( .A(B[30]), .B(B[31]), .Q(n149) );
  NOR24 U138 ( .A(net715654), .B(B[17]), .Q(n27) );
  NOR23 U139 ( .A(n66), .B(B[13]), .Q(n42) );
endmodule


module sqroot_comb_NBITS32_DW_cmp_47 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n28, n45, n47, n49, n51, n55, n57, n59, n85, net715492, net715628,
         net715660, net715592, n9, n82, n80, n8, n77, n76, n75, n74, n73, n72,
         n71, n70, n7, n69, n68, n67, n66, n65, n64, n63, n62, n61, n60, n6,
         n58, n56, n54, n52, n50, n5, n48, n46, n44, n43, n42, n41, n40, n4,
         n39, n38, n37, n36, n34, n32, n30, n3, n24, n22, n21, n20, n2, n19,
         n18, n17, n16, n15, n14, n13, n12, n11, n10, n1, n35, n33, n31, n29,
         n27, n26, n25, n23, n164, n165, n166, n167, n168, n169, n170, n171;

  NOR24 U2 ( .A(B[31]), .B(n2), .Q(n1) );
  OAI212 U41 ( .A(n41), .B(n52), .C(n42), .Q(n40) );
  OAI212 U63 ( .A(n66), .B(n63), .C(n64), .Q(n62) );
  AOI212 U39 ( .A(n39), .B(n62), .C(n40), .Q(n38) );
  OAI212 U70 ( .A(n70), .B(n73), .C(n71), .Q(n69) );
  OAI212 U75 ( .A(n77), .B(n75), .C(n76), .Q(n74) );
  AOI212 U68 ( .A(n74), .B(n68), .C(n69), .Q(n67) );
  OAI212 U37 ( .A(n37), .B(n67), .C(n38), .Q(n36) );
  AOI212 U12 ( .A(n36), .B(n12), .C(n13), .Q(n11) );
  NAND28 U1 ( .A(n11), .B(n1), .Q(GE_LT_GT_LE) );
  OAI212 U14 ( .A(n20), .B(n23), .C(n14), .Q(n13) );
  OAI212 U32 ( .A(n35), .B(n32), .C(n33), .Q(n31) );
  AOI212 U24 ( .A(n24), .B(n31), .C(n25), .Q(n23) );
  INV12 U97 ( .A(n45), .Q(n43) );
  NAND22 U98 ( .A(B[7]), .B(n168), .Q(n66) );
  NAND24 U99 ( .A(n19), .B(n21), .Q(n18) );
  INV3 U100 ( .A(n50), .Q(n48) );
  NOR24 U101 ( .A(n20), .B(n22), .Q(n12) );
  NAND21 U102 ( .A(B[5]), .B(n166), .Q(n73) );
  NAND22 U103 ( .A(B[14]), .B(n165), .Q(n33) );
  NAND26 U104 ( .A(n4), .B(n3), .Q(n2) );
  NOR24 U105 ( .A(n26), .B(n28), .Q(n24) );
  NAND22 U106 ( .A(B[13]), .B(net715592), .Q(n35) );
  INV3 U107 ( .A(A[13]), .Q(net715592) );
  NOR24 U108 ( .A(n165), .B(B[14]), .Q(n32) );
  INV3 U109 ( .A(A[14]), .Q(n165) );
  OAI212 U110 ( .A(n26), .B(n29), .C(n27), .Q(n25) );
  NOR24 U111 ( .A(n164), .B(B[16]), .Q(n26) );
  NAND26 U112 ( .A(B[15]), .B(net715660), .Q(n29) );
  INV3 U113 ( .A(A[15]), .Q(net715660) );
  NAND22 U114 ( .A(B[16]), .B(n164), .Q(n27) );
  INV3 U115 ( .A(A[16]), .Q(n164) );
  NAND23 U116 ( .A(n39), .B(n61), .Q(n37) );
  NOR24 U117 ( .A(n51), .B(n41), .Q(n39) );
  NOR22 U118 ( .A(n63), .B(n65), .Q(n61) );
  NOR24 U119 ( .A(n82), .B(B[8]), .Q(n63) );
  NOR22 U120 ( .A(n168), .B(B[7]), .Q(n65) );
  INV3 U121 ( .A(A[7]), .Q(n168) );
  NOR21 U122 ( .A(B[2]), .B(B[3]), .Q(n77) );
  NOR21 U123 ( .A(n167), .B(B[4]), .Q(n75) );
  INV1 U124 ( .A(A[4]), .Q(n167) );
  NAND20 U125 ( .A(B[4]), .B(n167), .Q(n76) );
  NOR22 U126 ( .A(n70), .B(n72), .Q(n68) );
  NOR24 U127 ( .A(n80), .B(B[6]), .Q(n70) );
  NOR21 U128 ( .A(n166), .B(B[5]), .Q(n72) );
  INV3 U129 ( .A(A[5]), .Q(n166) );
  NAND21 U130 ( .A(B[6]), .B(n80), .Q(n71) );
  INV0 U131 ( .A(A[6]), .Q(n80) );
  NAND21 U132 ( .A(B[8]), .B(n82), .Q(n64) );
  INV0 U133 ( .A(A[8]), .Q(n82) );
  NAND28 U134 ( .A(n47), .B(n43), .Q(n41) );
  AOI212 U135 ( .A(n58), .B(n171), .C(n54), .Q(n52) );
  CLKIN6 U136 ( .A(n60), .Q(n58) );
  NAND26 U137 ( .A(B[9]), .B(net715628), .Q(n60) );
  INV0 U138 ( .A(A[9]), .Q(net715628) );
  CLKIN6 U139 ( .A(n55), .Q(n171) );
  NOR24 U140 ( .A(n170), .B(B[10]), .Q(n55) );
  CLKIN4 U141 ( .A(n56), .Q(n54) );
  NAND22 U142 ( .A(B[10]), .B(n170), .Q(n56) );
  INV3 U143 ( .A(A[10]), .Q(n170) );
  AOI212 U144 ( .A(n43), .B(n48), .C(n44), .Q(n42) );
  NAND23 U145 ( .A(B[11]), .B(n85), .Q(n50) );
  INV3 U146 ( .A(A[11]), .Q(n85) );
  INV3 U147 ( .A(n46), .Q(n44) );
  NAND22 U148 ( .A(B[12]), .B(net715492), .Q(n46) );
  INV3 U149 ( .A(A[12]), .Q(net715492) );
  NOR24 U150 ( .A(n169), .B(B[17]), .Q(n20) );
  NAND23 U151 ( .A(n24), .B(n30), .Q(n22) );
  NOR22 U152 ( .A(n34), .B(n32), .Q(n30) );
  NOR24 U153 ( .A(net715592), .B(B[13]), .Q(n34) );
  NOR24 U154 ( .A(n18), .B(n15), .Q(n14) );
  NOR24 U155 ( .A(B[18]), .B(B[19]), .Q(n19) );
  NAND28 U156 ( .A(B[17]), .B(n169), .Q(n21) );
  INV3 U157 ( .A(A[17]), .Q(n169) );
  NAND24 U158 ( .A(n16), .B(n17), .Q(n15) );
  NOR24 U159 ( .A(B[23]), .B(B[22]), .Q(n16) );
  NOR23 U160 ( .A(B[21]), .B(B[20]), .Q(n17) );
  NOR24 U161 ( .A(n5), .B(n8), .Q(n4) );
  NAND24 U162 ( .A(n7), .B(n6), .Q(n5) );
  INV3 U163 ( .A(B[28]), .Q(n7) );
  INV6 U164 ( .A(B[29]), .Q(n6) );
  NAND24 U165 ( .A(n9), .B(n10), .Q(n8) );
  NOR24 U166 ( .A(B[26]), .B(B[27]), .Q(n9) );
  NOR24 U167 ( .A(B[25]), .B(B[24]), .Q(n10) );
  INV6 U168 ( .A(B[30]), .Q(n3) );
  INV6 U169 ( .A(n59), .Q(n57) );
  CLKIN6 U170 ( .A(n49), .Q(n47) );
  NAND24 U171 ( .A(n171), .B(n57), .Q(n51) );
  NOR24 U172 ( .A(net715660), .B(B[15]), .Q(n28) );
  NOR23 U173 ( .A(net715628), .B(B[9]), .Q(n59) );
  NOR24 U174 ( .A(n85), .B(B[11]), .Q(n49) );
  NOR24 U175 ( .A(net715492), .B(B[12]), .Q(n45) );
endmodule


module sqroot_comb_NBITS32_DW_cmp_49 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n66, n68, n71, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157;

  NOR24 U2 ( .A(B[31]), .B(n2), .Q(n1) );
  AOI212 U12 ( .A(n39), .B(n12), .C(n13), .Q(n11) );
  OAI212 U14 ( .A(n14), .B(n26), .C(n15), .Q(n13) );
  OAI212 U21 ( .A(n21), .B(n24), .C(n22), .Q(n20) );
  AOI212 U27 ( .A(n27), .B(n34), .C(n28), .Q(n26) );
  OAI212 U29 ( .A(n32), .B(n29), .C(n30), .Q(n28) );
  NOR24 U30 ( .A(n148), .B(B[16]), .Q(n29) );
  OAI212 U35 ( .A(n38), .B(n35), .C(n36), .Q(n34) );
  OAI212 U40 ( .A(n40), .B(n54), .C(n41), .Q(n39) );
  AOI212 U55 ( .A(n61), .B(n55), .C(n56), .Q(n54) );
  NOR23 U83 ( .A(B[26]), .B(B[25]), .Q(n9) );
  NAND21 U84 ( .A(B[12]), .B(n71), .Q(n45) );
  NOR24 U85 ( .A(n149), .B(B[10]), .Q(n50) );
  NOR24 U86 ( .A(B[24]), .B(B[23]), .Q(n10) );
  NAND23 U87 ( .A(B[13]), .B(n153), .Q(n38) );
  NAND26 U88 ( .A(n4), .B(n3), .Q(n2) );
  NAND28 U89 ( .A(n18), .B(n17), .Q(n16) );
  NOR22 U90 ( .A(n157), .B(B[6]), .Q(n62) );
  OAI212 U91 ( .A(n62), .B(n64), .C(n63), .Q(n61) );
  NAND26 U92 ( .A(n11), .B(n1), .Q(GE_LT_GT_LE) );
  NOR24 U93 ( .A(n156), .B(B[8]), .Q(n57) );
  NOR23 U94 ( .A(n59), .B(n57), .Q(n55) );
  OAI212 U95 ( .A(n60), .B(n57), .C(n58), .Q(n56) );
  NOR22 U96 ( .A(n66), .B(B[7]), .Q(n59) );
  NOR23 U97 ( .A(n37), .B(n35), .Q(n33) );
  NOR22 U98 ( .A(B[4]), .B(B[5]), .Q(n64) );
  NOR23 U99 ( .A(n16), .B(n20), .Q(n15) );
  NOR23 U100 ( .A(n151), .B(B[15]), .Q(n31) );
  OAI212 U101 ( .A(n44), .B(n47), .C(n45), .Q(n43) );
  CLKIN2 U102 ( .A(A[6]), .Q(n157) );
  NOR24 U103 ( .A(n21), .B(n23), .Q(n19) );
  NAND26 U104 ( .A(n7), .B(n6), .Q(n5) );
  NOR23 U105 ( .A(B[28]), .B(B[27]), .Q(n7) );
  NAND24 U106 ( .A(n9), .B(n10), .Q(n8) );
  NOR23 U107 ( .A(n31), .B(n29), .Q(n27) );
  NAND23 U108 ( .A(B[17]), .B(n154), .Q(n24) );
  NAND23 U109 ( .A(B[15]), .B(n151), .Q(n32) );
  NOR23 U110 ( .A(n154), .B(B[17]), .Q(n23) );
  NAND24 U111 ( .A(n27), .B(n33), .Q(n25) );
  NOR24 U112 ( .A(n5), .B(n8), .Q(n4) );
  CLKIN3 U113 ( .A(A[10]), .Q(n149) );
  NOR23 U114 ( .A(n150), .B(B[14]), .Q(n35) );
  NOR22 U115 ( .A(n152), .B(B[11]), .Q(n46) );
  NOR23 U116 ( .A(n14), .B(n25), .Q(n12) );
  NOR23 U117 ( .A(n153), .B(B[13]), .Q(n37) );
  NAND22 U118 ( .A(B[11]), .B(n152), .Q(n47) );
  NOR24 U119 ( .A(B[20]), .B(B[19]), .Q(n18) );
  NOR24 U120 ( .A(B[22]), .B(B[21]), .Q(n17) );
  NOR22 U121 ( .A(n68), .B(B[9]), .Q(n52) );
  INV6 U122 ( .A(n19), .Q(n14) );
  NOR22 U123 ( .A(n50), .B(n52), .Q(n48) );
  OAI211 U124 ( .A(n53), .B(n50), .C(n51), .Q(n49) );
  NAND22 U125 ( .A(B[9]), .B(n68), .Q(n53) );
  NAND21 U126 ( .A(B[10]), .B(n149), .Q(n51) );
  NAND21 U127 ( .A(B[8]), .B(n156), .Q(n58) );
  NOR23 U128 ( .A(n71), .B(B[12]), .Q(n44) );
  NOR23 U129 ( .A(n46), .B(n44), .Q(n42) );
  NOR24 U130 ( .A(n155), .B(B[18]), .Q(n21) );
  NAND21 U131 ( .A(B[18]), .B(n155), .Q(n22) );
  NAND22 U132 ( .A(B[7]), .B(n66), .Q(n60) );
  INV0 U133 ( .A(A[9]), .Q(n68) );
  NAND21 U134 ( .A(B[14]), .B(n150), .Q(n36) );
  AOI212 U135 ( .A(n49), .B(n42), .C(n43), .Q(n41) );
  NAND21 U136 ( .A(B[6]), .B(n157), .Q(n63) );
  INV6 U137 ( .A(B[30]), .Q(n3) );
  CLKIN0 U138 ( .A(A[11]), .Q(n152) );
  INV0 U139 ( .A(A[12]), .Q(n71) );
  CLKIN0 U140 ( .A(A[7]), .Q(n66) );
  INV3 U141 ( .A(A[8]), .Q(n156) );
  INV3 U142 ( .A(B[29]), .Q(n6) );
  INV3 U143 ( .A(A[13]), .Q(n153) );
  INV3 U144 ( .A(A[14]), .Q(n150) );
  INV3 U145 ( .A(A[15]), .Q(n151) );
  INV3 U146 ( .A(A[17]), .Q(n154) );
  INV3 U147 ( .A(A[16]), .Q(n148) );
  INV3 U148 ( .A(A[18]), .Q(n155) );
  NAND22 U149 ( .A(n48), .B(n42), .Q(n40) );
  NAND21 U150 ( .A(B[16]), .B(n148), .Q(n30) );
endmodule


module sqroot_comb_NBITS32_DW_cmp_50 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n22, n30, n32, n34, n57, n59, n61, n69, n104, net715434, net715468,
         net715528, net715632, net715664, net719411, net722375, net722374,
         net715596, n99, n95, n94, n93, n92, n91, n90, n9, n89, n88, n87, n86,
         n85, n84, n83, n82, n81, n80, n8, n78, n76, n75, n74, n72, n70, n7,
         n68, n67, n66, n65, n64, n63, n62, n60, n6, n58, n56, n54, n52, n51,
         n50, n5, n49, n48, n47, n46, n44, n42, n4, n36, n3, n26, n24, n2, n17,
         n15, n14, n13, n12, n11, n101, n10, n1, n35, n33, n31, n29, n28, n27,
         n25, n23, n21, n20, n19, n18, n16, net715560, n45, n43, n41, n40, n39,
         n38, n37, n185, n186, n187, n188, n189, n190, n191, n192, n193;

  OAI212 U51 ( .A(n62), .B(n51), .C(n52), .Q(n50) );
  AOI212 U77 ( .A(n193), .B(n82), .C(n78), .Q(n76) );
  OAI212 U65 ( .A(n65), .B(n76), .C(n66), .Q(n64) );
  OAI212 U88 ( .A(n91), .B(n88), .C(n89), .Q(n87) );
  OAI212 U93 ( .A(n93), .B(n95), .C(n94), .Q(n92) );
  AOI212 U86 ( .A(n92), .B(n86), .C(n87), .Q(n85) );
  OAI212 U47 ( .A(n47), .B(n85), .C(n48), .Q(n46) );
  AOI212 U6 ( .A(n46), .B(n6), .C(n7), .Q(n5) );
  AOI212 U17 ( .A(n25), .B(n17), .C(n18), .Q(n16) );
  OAI212 U26 ( .A(n26), .B(n37), .C(n27), .Q(n25) );
  NAND24 U116 ( .A(n24), .B(n17), .Q(n15) );
  NAND23 U117 ( .A(B[14]), .B(net715664), .Q(n35) );
  CLKIN6 U118 ( .A(B[6]), .Q(n191) );
  NAND22 U119 ( .A(B[6]), .B(n188), .Q(n80) );
  NOR23 U120 ( .A(n36), .B(n26), .Q(n24) );
  NOR22 U121 ( .A(n186), .B(B[3]), .Q(n90) );
  NOR23 U122 ( .A(n185), .B(B[4]), .Q(n88) );
  INV6 U123 ( .A(n45), .Q(n43) );
  INV10 U124 ( .A(B[7]), .Q(net722375) );
  NAND28 U125 ( .A(n191), .B(n190), .Q(n193) );
  INV6 U126 ( .A(n35), .Q(n33) );
  NOR24 U127 ( .A(n90), .B(n88), .Q(n86) );
  INV8 U128 ( .A(n69), .Q(n67) );
  NAND21 U129 ( .A(B[4]), .B(n185), .Q(n89) );
  CLKIN3 U130 ( .A(n56), .Q(n54) );
  CLKIN12 U131 ( .A(B[11]), .Q(net719411) );
  INV3 U132 ( .A(n188), .Q(n190) );
  AOI212 U133 ( .A(n38), .B(n43), .C(n39), .Q(n37) );
  INV6 U134 ( .A(n40), .Q(n38) );
  NAND28 U135 ( .A(B[12]), .B(net715596), .Q(n45) );
  INV3 U136 ( .A(A[12]), .Q(net715596) );
  INV4 U137 ( .A(n41), .Q(n39) );
  NAND23 U138 ( .A(B[13]), .B(net715560), .Q(n41) );
  INV3 U139 ( .A(A[13]), .Q(net715560) );
  NOR24 U140 ( .A(net715560), .B(B[13]), .Q(n40) );
  NAND22 U141 ( .A(n38), .B(n42), .Q(n36) );
  NAND24 U142 ( .A(n32), .B(n28), .Q(n26) );
  AOI212 U143 ( .A(n28), .B(n33), .C(n29), .Q(n27) );
  INV6 U144 ( .A(n30), .Q(n28) );
  INV3 U145 ( .A(A[14]), .Q(net715664) );
  INV3 U146 ( .A(n31), .Q(n29) );
  NAND22 U147 ( .A(B[15]), .B(net715468), .Q(n31) );
  INV1 U148 ( .A(A[15]), .Q(net715468) );
  INV6 U149 ( .A(n22), .Q(n17) );
  NAND24 U150 ( .A(n19), .B(n20), .Q(n18) );
  NOR23 U151 ( .A(B[19]), .B(B[18]), .Q(n19) );
  NOR24 U152 ( .A(n21), .B(B[17]), .Q(n20) );
  CLKIN6 U153 ( .A(n23), .Q(n21) );
  NAND26 U154 ( .A(B[16]), .B(net715434), .Q(n23) );
  INV3 U155 ( .A(A[16]), .Q(net715434) );
  NAND24 U156 ( .A(n8), .B(n16), .Q(n7) );
  NAND26 U157 ( .A(n5), .B(n1), .Q(GE_LT_GT_LE) );
  NAND24 U158 ( .A(n49), .B(n63), .Q(n47) );
  NOR24 U159 ( .A(n61), .B(n51), .Q(n49) );
  NOR24 U160 ( .A(n65), .B(n75), .Q(n63) );
  NAND28 U161 ( .A(n67), .B(net722374), .Q(n65) );
  NAND24 U162 ( .A(n81), .B(n193), .Q(n75) );
  INV2 U163 ( .A(n83), .Q(n81) );
  NOR21 U164 ( .A(n99), .B(B[5]), .Q(n83) );
  INV0 U165 ( .A(A[5]), .Q(n99) );
  NOR23 U166 ( .A(n187), .B(B[2]), .Q(n93) );
  INV1 U167 ( .A(A[2]), .Q(n187) );
  NOR24 U168 ( .A(B[1]), .B(B[0]), .Q(n95) );
  NAND21 U169 ( .A(B[2]), .B(n187), .Q(n94) );
  INV0 U170 ( .A(A[3]), .Q(n186) );
  NAND21 U171 ( .A(B[3]), .B(n186), .Q(n91) );
  INV3 U172 ( .A(A[4]), .Q(n185) );
  AOI212 U173 ( .A(n64), .B(n49), .C(n50), .Q(n48) );
  INV3 U174 ( .A(n84), .Q(n82) );
  NAND22 U175 ( .A(B[5]), .B(n99), .Q(n84) );
  INV3 U176 ( .A(n80), .Q(n78) );
  INV3 U177 ( .A(A[6]), .Q(n188) );
  AOI212 U178 ( .A(n67), .B(n72), .C(n68), .Q(n66) );
  INV6 U179 ( .A(n74), .Q(n72) );
  NAND24 U180 ( .A(B[7]), .B(n101), .Q(n74) );
  INV0 U181 ( .A(A[7]), .Q(n101) );
  INV3 U182 ( .A(n70), .Q(n68) );
  NAND22 U183 ( .A(B[8]), .B(net715632), .Q(n70) );
  INV3 U184 ( .A(A[8]), .Q(net715632) );
  NAND22 U185 ( .A(B[9]), .B(net715528), .Q(n62) );
  INV3 U186 ( .A(A[9]), .Q(net715528) );
  NAND28 U187 ( .A(n57), .B(n192), .Q(n51) );
  AOI212 U188 ( .A(n58), .B(n192), .C(n54), .Q(n52) );
  INV2 U189 ( .A(n60), .Q(n58) );
  NAND22 U190 ( .A(B[10]), .B(n104), .Q(n60) );
  INV3 U191 ( .A(A[10]), .Q(n104) );
  NAND28 U192 ( .A(net719411), .B(A[11]), .Q(n192) );
  NAND22 U193 ( .A(B[11]), .B(n189), .Q(n56) );
  INV0 U194 ( .A(A[11]), .Q(n189) );
  INV6 U195 ( .A(n15), .Q(n6) );
  INV3 U196 ( .A(n44), .Q(n42) );
  NOR24 U197 ( .A(net715596), .B(B[12]), .Q(n44) );
  NOR24 U198 ( .A(n12), .B(n9), .Q(n8) );
  NAND24 U199 ( .A(n14), .B(n13), .Q(n12) );
  NOR24 U200 ( .A(B[20]), .B(B[21]), .Q(n14) );
  NOR24 U201 ( .A(B[23]), .B(B[22]), .Q(n13) );
  NAND24 U202 ( .A(n10), .B(n11), .Q(n9) );
  NOR24 U203 ( .A(B[26]), .B(B[27]), .Q(n10) );
  NOR23 U204 ( .A(B[24]), .B(B[25]), .Q(n11) );
  NOR24 U205 ( .A(B[31]), .B(n2), .Q(n1) );
  NAND24 U206 ( .A(n4), .B(n3), .Q(n2) );
  NOR23 U207 ( .A(B[29]), .B(B[28]), .Q(n4) );
  INV3 U208 ( .A(B[30]), .Q(n3) );
  NAND28 U209 ( .A(A[7]), .B(net722375), .Q(net722374) );
  NOR23 U210 ( .A(n104), .B(B[10]), .Q(n59) );
  CLKIN6 U211 ( .A(n34), .Q(n32) );
  NOR24 U212 ( .A(net715468), .B(B[15]), .Q(n30) );
  NOR23 U213 ( .A(net715528), .B(B[9]), .Q(n61) );
  NOR24 U214 ( .A(net715664), .B(B[14]), .Q(n34) );
  NOR24 U215 ( .A(net715434), .B(B[16]), .Q(n22) );
  NOR24 U216 ( .A(net715632), .B(B[8]), .Q(n69) );
  INV3 U217 ( .A(n59), .Q(n57) );
endmodule


module sqroot_comb_NBITS32_DW01_sub_69 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n14, n15, n16, n18, n19, n20, n21, n22, n23, n24, n25, n26, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n42, n43, n46,
         n47, n48, n51, n54, n55, n58, n59, n60, n64, n65, n69, n70, n73, n74,
         n77, n78, n79, n81, n82, n85, n86, n87, n89, n90, n91, n95, n97, n98,
         n99, n100, n103, n105, n107, n109, n112, n113, n114, n115, n116, n118,
         n119, n120, n121, n122, n123, n124, n125, n128, n129, n130, n131,
         n132, n133, n134, n136, n137, n138, n141, n142, n143, n148, n149,
         n150, n151, n152, n153, n160, n161, n162, n163, n164, n167, n168,
         n169, n170, n171, n172, n175, n176, n177, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n220, n222, net715530, net715562, net715848,
         net718538, net718537, net723451, n17, n140, n139, n157, n156, n155,
         n154, n217, n159, n158, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344;

  OAI212 U111 ( .A(n120), .B(n112), .C(n113), .Q(n107) );
  NOR24 U124 ( .A(n341), .B(A[17]), .Q(n119) );
  AOI212 U133 ( .A(n128), .B(n143), .C(n129), .Q(n123) );
  OAI212 U135 ( .A(n138), .B(n130), .C(n131), .Q(n129) );
  OAI212 U141 ( .A(n153), .B(n133), .C(n134), .Q(n132) );
  OAI212 U215 ( .A(n190), .B(n186), .C(n187), .Q(n185) );
  OAI212 U228 ( .A(n193), .B(n195), .C(n194), .Q(n192) );
  OAI212 U151 ( .A(n153), .B(n140), .C(n141), .Q(n139) );
  AOI212 U60 ( .A(n154), .B(n69), .C(n70), .Q(n1) );
  OAI212 U198 ( .A(n181), .B(n175), .C(n176), .Q(n170) );
  AOI212 U213 ( .A(n184), .B(n192), .C(n185), .Q(n183) );
  OAI212 U172 ( .A(n183), .B(n155), .C(n156), .Q(n154) );
  AOI212 U174 ( .A(n157), .B(n170), .C(n158), .Q(n156) );
  OAI212 U176 ( .A(n159), .B(n167), .C(n160), .Q(n158) );
  INV3 U255 ( .A(n90), .Q(n91) );
  INV3 U256 ( .A(n170), .Q(n172) );
  INV2 U257 ( .A(n125), .Q(n327) );
  NOR23 U258 ( .A(n337), .B(A[16]), .Q(n130) );
  INV3 U259 ( .A(net718537), .Q(n318) );
  INV2 U260 ( .A(B[6]), .Q(n344) );
  XOR20 U261 ( .A(n19), .B(n153), .Q(DIFF[13]) );
  INV1 U262 ( .A(n137), .Q(n201) );
  NOR22 U263 ( .A(n34), .B(n48), .Q(n33) );
  NAND22 U264 ( .A(n332), .B(n333), .Q(DIFF[28]) );
  NAND22 U265 ( .A(A[14]), .B(n339), .Q(n149) );
  INV0 U266 ( .A(n143), .Q(n141) );
  NAND22 U267 ( .A(n124), .B(n98), .Q(n78) );
  INV6 U268 ( .A(n107), .Q(n109) );
  INV0 U269 ( .A(n175), .Q(n206) );
  NOR24 U270 ( .A(net715562), .B(A[15]), .Q(n137) );
  NOR22 U271 ( .A(A[4]), .B(A[5]), .Q(n319) );
  INV3 U272 ( .A(n20), .Q(n329) );
  NOR24 U273 ( .A(n217), .B(A[12]), .Q(n159) );
  NAND26 U274 ( .A(A[11]), .B(net715530), .Q(n167) );
  NAND22 U275 ( .A(A[12]), .B(n217), .Q(n160) );
  INV0 U276 ( .A(B[12]), .Q(n217) );
  NOR22 U277 ( .A(n159), .B(n164), .Q(n157) );
  INV0 U278 ( .A(n159), .Q(n204) );
  NAND22 U279 ( .A(n157), .B(n169), .Q(n155) );
  NOR24 U280 ( .A(n175), .B(n180), .Q(n169) );
  INV8 U281 ( .A(n154), .Q(n153) );
  XNR22 U282 ( .A(n17), .B(n139), .Q(DIFF[15]) );
  NAND21 U283 ( .A(n201), .B(n138), .Q(n17) );
  NAND22 U284 ( .A(A[15]), .B(net715562), .Q(n138) );
  INV3 U285 ( .A(n142), .Q(n140) );
  NOR23 U286 ( .A(n148), .B(n151), .Q(n142) );
  NOR23 U287 ( .A(n189), .B(n325), .Q(n184) );
  INV1 U288 ( .A(n112), .Q(n198) );
  XNR22 U289 ( .A(n85), .B(A[21]), .Q(DIFF[21]) );
  NAND22 U290 ( .A(n15), .B(n335), .Q(n322) );
  NAND24 U291 ( .A(n320), .B(n321), .Q(n323) );
  NAND24 U292 ( .A(n322), .B(n323), .Q(DIFF[17]) );
  INV2 U293 ( .A(n15), .Q(n320) );
  CLKIN6 U294 ( .A(n335), .Q(n321) );
  NAND22 U295 ( .A(n199), .B(n120), .Q(n15) );
  OAI211 U296 ( .A(n172), .B(n164), .C(n167), .Q(n163) );
  NOR21 U297 ( .A(A[22]), .B(A[21]), .Q(n74) );
  CLKIN1 U298 ( .A(A[23]), .Q(n65) );
  CLKIN3 U299 ( .A(n172), .Q(net723451) );
  XOR21 U300 ( .A(n25), .B(n191), .Q(DIFF[7]) );
  INV2 U301 ( .A(A[19]), .Q(n100) );
  NAND21 U302 ( .A(n187), .B(n208), .Q(n24) );
  NOR23 U303 ( .A(n343), .B(A[8]), .Q(n186) );
  NAND24 U304 ( .A(A[6]), .B(n344), .Q(n194) );
  AOI211 U305 ( .A(n125), .B(n199), .C(n118), .Q(n116) );
  OAI2112 U306 ( .A(n336), .B(n123), .C(n324), .D(n109), .Q(n70) );
  INV3 U307 ( .A(n73), .Q(n324) );
  NAND21 U308 ( .A(net715848), .B(n33), .Q(n32) );
  NOR23 U309 ( .A(n343), .B(A[8]), .Q(n325) );
  OAI212 U310 ( .A(n78), .B(n153), .C(n97), .Q(n95) );
  INV0 U311 ( .A(n325), .Q(n208) );
  OAI210 U312 ( .A(n193), .B(n319), .C(n194), .Q(n326) );
  NAND23 U313 ( .A(net715848), .B(n43), .Q(n42) );
  XNR21 U314 ( .A(A[27]), .B(n46), .Q(DIFF[27]) );
  XNR21 U315 ( .A(A[30]), .B(n32), .Q(DIFF[30]) );
  NOR24 U316 ( .A(n137), .B(n130), .Q(n128) );
  XNR20 U317 ( .A(A[4]), .B(A[5]), .Q(DIFF[5]) );
  NAND24 U318 ( .A(A[17]), .B(n341), .Q(n120) );
  NAND22 U319 ( .A(n124), .B(n199), .Q(n115) );
  INV1 U320 ( .A(n119), .Q(n199) );
  NAND23 U321 ( .A(net715848), .B(n59), .Q(n58) );
  NAND23 U322 ( .A(net715848), .B(n37), .Q(n36) );
  NAND23 U323 ( .A(net715848), .B(n65), .Q(n64) );
  NAND23 U324 ( .A(net715848), .B(n55), .Q(n54) );
  INV1 U325 ( .A(n326), .Q(n191) );
  NAND26 U326 ( .A(A[9]), .B(n220), .Q(n181) );
  NOR23 U327 ( .A(n220), .B(A[9]), .Q(n180) );
  CLKBU15 U328 ( .A(n1), .Q(net715848) );
  INV6 U329 ( .A(n123), .Q(n125) );
  NAND20 U330 ( .A(n205), .B(n167), .Q(n21) );
  NOR24 U331 ( .A(n222), .B(A[7]), .Q(n189) );
  CLKIN12 U332 ( .A(n98), .Q(n336) );
  BUF2 U333 ( .A(n319), .Q(n328) );
  NAND22 U334 ( .A(n210), .B(n194), .Q(n26) );
  CLKIN0 U335 ( .A(n130), .Q(n200) );
  XNR21 U336 ( .A(n23), .B(n318), .Q(DIFF[9]) );
  AOI212 U337 ( .A(n125), .B(n98), .C(n89), .Q(n87) );
  NOR23 U338 ( .A(net723451), .B(n334), .Q(n168) );
  XNR22 U339 ( .A(n24), .B(n188), .Q(DIFF[8]) );
  NAND21 U340 ( .A(A[18]), .B(n342), .Q(n113) );
  XOR22 U341 ( .A(A[23]), .B(net715848), .Q(DIFF[23]) );
  NOR22 U342 ( .A(n336), .B(n122), .Q(n69) );
  NOR24 U343 ( .A(A[20]), .B(A[19]), .Q(n90) );
  NOR24 U344 ( .A(net718537), .B(net718538), .Q(n334) );
  NAND23 U345 ( .A(net715848), .B(n47), .Q(n46) );
  CLKIN6 U346 ( .A(n182), .Q(net718537) );
  NOR24 U347 ( .A(n344), .B(A[6]), .Q(n193) );
  NOR21 U348 ( .A(A[28]), .B(A[27]), .Q(n39) );
  NAND22 U349 ( .A(A[8]), .B(n343), .Q(n187) );
  OAI210 U350 ( .A(n153), .B(n122), .C(n327), .Q(n121) );
  NAND22 U351 ( .A(A[16]), .B(n337), .Q(n131) );
  INV1 U352 ( .A(n39), .Q(n38) );
  NAND21 U353 ( .A(n124), .B(n98), .Q(n86) );
  XOR22 U354 ( .A(n22), .B(n177), .Q(DIFF[10]) );
  OAI212 U355 ( .A(n153), .B(n86), .C(n87), .Q(n85) );
  XNR22 U356 ( .A(A[24]), .B(n64), .Q(DIFF[24]) );
  OAI211 U357 ( .A(n115), .B(n153), .C(n116), .Q(n114) );
  OAI211 U358 ( .A(n78), .B(n153), .C(n79), .Q(n77) );
  OAI211 U359 ( .A(n153), .B(n78), .C(n105), .Q(n103) );
  NOR21 U360 ( .A(n38), .B(n48), .Q(n37) );
  INV4 U361 ( .A(n183), .Q(n182) );
  XNR22 U362 ( .A(A[25]), .B(n58), .Q(DIFF[25]) );
  XNR22 U363 ( .A(n329), .B(n161), .Q(DIFF[12]) );
  INV6 U364 ( .A(n122), .Q(n124) );
  XNR21 U365 ( .A(A[22]), .B(n77), .Q(DIFF[22]) );
  NAND21 U366 ( .A(net715848), .B(n29), .Q(n28) );
  NAND21 U367 ( .A(n33), .B(n31), .Q(n30) );
  NAND21 U368 ( .A(A[28]), .B(n42), .Q(n332) );
  CLKIN0 U369 ( .A(A[28]), .Q(n330) );
  NAND22 U370 ( .A(n109), .B(n90), .Q(n89) );
  AOI211 U371 ( .A(n125), .B(n98), .C(n107), .Q(n105) );
  XNR22 U372 ( .A(n14), .B(n114), .Q(DIFF[18]) );
  OAI211 U373 ( .A(n189), .B(n191), .C(n190), .Q(n188) );
  XNR21 U374 ( .A(A[20]), .B(n95), .Q(DIFF[20]) );
  NOR24 U375 ( .A(n340), .B(A[13]), .Q(n151) );
  XNR22 U376 ( .A(n18), .B(n150), .Q(DIFF[14]) );
  NAND21 U377 ( .A(n200), .B(n131), .Q(n16) );
  XNR22 U378 ( .A(n16), .B(n132), .Q(DIFF[16]) );
  XNR22 U379 ( .A(A[26]), .B(n54), .Q(DIFF[26]) );
  AOI212 U380 ( .A(n182), .B(n207), .C(n179), .Q(n177) );
  CLKIN0 U381 ( .A(B[7]), .Q(n222) );
  OAI212 U382 ( .A(n153), .B(n151), .C(n152), .Q(n150) );
  NOR24 U383 ( .A(n339), .B(A[14]), .Q(n148) );
  XNR22 U384 ( .A(A[29]), .B(n36), .Q(DIFF[29]) );
  NOR24 U385 ( .A(n338), .B(A[10]), .Q(n175) );
  NAND21 U386 ( .A(n109), .B(n82), .Q(n81) );
  NAND22 U387 ( .A(n109), .B(n100), .Q(n99) );
  NOR24 U388 ( .A(net715530), .B(A[11]), .Q(n164) );
  NOR24 U389 ( .A(n112), .B(n119), .Q(n98) );
  NAND22 U390 ( .A(n330), .B(n331), .Q(n333) );
  CLKIN3 U391 ( .A(n42), .Q(n331) );
  INV1 U392 ( .A(n169), .Q(net718538) );
  XOR22 U393 ( .A(n21), .B(n168), .Q(DIFF[11]) );
  XNR21 U394 ( .A(A[31]), .B(n28), .Q(DIFF[31]) );
  AOI211 U395 ( .A(n125), .B(n98), .C(n99), .Q(n97) );
  AOI212 U396 ( .A(n182), .B(n162), .C(n163), .Q(n161) );
  XNR21 U397 ( .A(A[19]), .B(n103), .Q(DIFF[19]) );
  NAND22 U398 ( .A(n206), .B(n176), .Q(n22) );
  NAND22 U399 ( .A(A[10]), .B(n338), .Q(n176) );
  NOR24 U400 ( .A(A[4]), .B(A[5]), .Q(n195) );
  NOR24 U401 ( .A(n342), .B(A[18]), .Q(n112) );
  INV6 U402 ( .A(n180), .Q(n207) );
  NAND22 U403 ( .A(n203), .B(n152), .Q(n19) );
  OAI212 U404 ( .A(n152), .B(n148), .C(n149), .Q(n143) );
  NAND24 U405 ( .A(A[13]), .B(n340), .Q(n152) );
  CLKIN2 U406 ( .A(n59), .Q(n60) );
  NAND24 U407 ( .A(n51), .B(n59), .Q(n48) );
  NOR24 U408 ( .A(A[24]), .B(A[23]), .Q(n59) );
  NAND22 U409 ( .A(A[7]), .B(n222), .Q(n190) );
  INV3 U410 ( .A(n148), .Q(n202) );
  CLKIN3 U411 ( .A(n169), .Q(n171) );
  CLKIN0 U412 ( .A(n189), .Q(n209) );
  NAND20 U413 ( .A(n207), .B(n181), .Q(n23) );
  NAND24 U414 ( .A(n128), .B(n142), .Q(n122) );
  NAND20 U415 ( .A(n198), .B(n113), .Q(n14) );
  INV0 U416 ( .A(B[9]), .Q(n220) );
  INV0 U417 ( .A(n48), .Q(n47) );
  INV0 U418 ( .A(n151), .Q(n203) );
  INV0 U419 ( .A(B[10]), .Q(n338) );
  NOR20 U420 ( .A(A[21]), .B(n91), .Q(n82) );
  INV0 U421 ( .A(n164), .Q(n205) );
  NOR21 U422 ( .A(n164), .B(n171), .Q(n162) );
  INV0 U423 ( .A(n120), .Q(n118) );
  NAND21 U424 ( .A(n160), .B(n204), .Q(n20) );
  CLKIN0 U425 ( .A(B[11]), .Q(net715530) );
  INV0 U426 ( .A(n193), .Q(n210) );
  NAND20 U427 ( .A(n209), .B(n190), .Q(n25) );
  XOR20 U428 ( .A(n328), .B(n26), .Q(DIFF[6]) );
  INV3 U429 ( .A(B[8]), .Q(n343) );
  AOI211 U430 ( .A(n125), .B(n98), .C(n81), .Q(n79) );
  NAND22 U431 ( .A(n39), .B(n35), .Q(n34) );
  INV0 U432 ( .A(A[29]), .Q(n35) );
  NOR20 U433 ( .A(A[25]), .B(n60), .Q(n55) );
  INV3 U434 ( .A(n30), .Q(n29) );
  INV0 U435 ( .A(A[30]), .Q(n31) );
  NAND22 U436 ( .A(n202), .B(n149), .Q(n18) );
  NAND22 U437 ( .A(n142), .B(n201), .Q(n133) );
  AOI210 U438 ( .A(n143), .B(n201), .C(n136), .Q(n134) );
  INV3 U439 ( .A(n138), .Q(n136) );
  NAND22 U440 ( .A(n74), .B(n90), .Q(n73) );
  INV3 U441 ( .A(B[13]), .Q(n340) );
  INV3 U442 ( .A(B[14]), .Q(n339) );
  INV3 U443 ( .A(B[15]), .Q(net715562) );
  INV3 U444 ( .A(B[17]), .Q(n341) );
  INV3 U445 ( .A(n181), .Q(n179) );
  INV3 U446 ( .A(B[16]), .Q(n337) );
  INV3 U447 ( .A(B[18]), .Q(n342) );
  BUF6 U448 ( .A(n121), .Q(n335) );
  NOR21 U449 ( .A(A[27]), .B(n48), .Q(n43) );
  NOR21 U450 ( .A(A[26]), .B(A[25]), .Q(n51) );
endmodule


module sqroot_comb_NBITS32_DW_cmp_48 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n22, n24, n26, n30, n32, n34, n49, n59, n74, n76, n90, net715318,
         net715472, net715532, net715564, n93, n9, n8, n7, n64, n63, n62, n61,
         n6, n57, n56, n55, n54, n53, n52, n51, n50, n5, n48, n47, n46, n45,
         n44, n43, n42, n41, n40, n4, n39, n38, n37, n36, n35, n33, n31, n3,
         n29, n28, n27, n25, n23, n21, n20, n19, n18, n17, n16, n15, n14, n13,
         n12, n11, n10, n83, n82, n81, n80, n79, n78, n68, n67, n66, n65, n88,
         n77, n75, n73, n72, n71, n70, n69, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190;

  OAI212 U17 ( .A(n17), .B(n29), .C(n18), .Q(n16) );
  OAI212 U47 ( .A(n50), .B(n47), .C(n48), .Q(n46) );
  OAI212 U53 ( .A(n53), .B(n56), .C(n54), .Q(n52) );
  OAI212 U43 ( .A(n43), .B(n65), .C(n44), .Q(n42) );
  OAI212 U81 ( .A(n81), .B(n83), .C(n82), .Q(n80) );
  OAI212 U68 ( .A(n79), .B(n68), .C(n69), .Q(n67) );
  NAND23 U105 ( .A(n190), .B(n36), .Q(n28) );
  NAND23 U106 ( .A(B[2]), .B(n174), .Q(n79) );
  NAND24 U107 ( .A(n51), .B(n45), .Q(n43) );
  CLKIN6 U108 ( .A(n22), .Q(n17) );
  NOR24 U109 ( .A(B[16]), .B(B[17]), .Q(n21) );
  CLKIN1 U110 ( .A(A[0]), .Q(n176) );
  NAND23 U111 ( .A(n3), .B(n187), .Q(n186) );
  INV4 U112 ( .A(n37), .Q(n183) );
  NOR22 U113 ( .A(n177), .B(B[5]), .Q(n63) );
  NAND23 U114 ( .A(B[5]), .B(n177), .Q(n64) );
  NOR23 U115 ( .A(B[19]), .B(B[18]), .Q(n20) );
  INV3 U116 ( .A(B[31]), .Q(n187) );
  AOI212 U117 ( .A(n70), .B(n75), .C(n71), .Q(n69) );
  CLKIN6 U118 ( .A(n72), .Q(n70) );
  INV3 U119 ( .A(n77), .Q(n75) );
  NAND23 U120 ( .A(B[3]), .B(net715318), .Q(n77) );
  INV3 U121 ( .A(A[3]), .Q(net715318) );
  CLKIN3 U122 ( .A(n73), .Q(n71) );
  NAND21 U123 ( .A(B[4]), .B(n88), .Q(n73) );
  INV0 U124 ( .A(A[4]), .Q(n88) );
  NOR23 U125 ( .A(n88), .B(B[4]), .Q(n72) );
  NAND24 U126 ( .A(n74), .B(n70), .Q(n68) );
  AOI212 U127 ( .A(n66), .B(n80), .C(n67), .Q(n65) );
  NOR22 U128 ( .A(n78), .B(n68), .Q(n66) );
  NOR22 U129 ( .A(n174), .B(B[2]), .Q(n78) );
  CLKIN0 U130 ( .A(A[2]), .Q(n174) );
  NOR23 U131 ( .A(n175), .B(B[1]), .Q(n81) );
  INV0 U132 ( .A(A[1]), .Q(n175) );
  NAND22 U133 ( .A(B[0]), .B(n176), .Q(n83) );
  NAND21 U134 ( .A(B[1]), .B(n175), .Q(n82) );
  NAND24 U135 ( .A(n14), .B(n188), .Q(GE_LT_GT_LE) );
  AOI212 U136 ( .A(n42), .B(n15), .C(n16), .Q(n14) );
  NOR22 U137 ( .A(n53), .B(n55), .Q(n51) );
  NOR24 U138 ( .A(n181), .B(B[7]), .Q(n53) );
  NAND22 U139 ( .A(n57), .B(n61), .Q(n55) );
  CLKIN6 U140 ( .A(n59), .Q(n57) );
  INV3 U141 ( .A(n63), .Q(n61) );
  INV3 U142 ( .A(A[5]), .Q(n177) );
  NOR23 U143 ( .A(n49), .B(n47), .Q(n45) );
  AOI212 U144 ( .A(n52), .B(n45), .C(n46), .Q(n44) );
  AOI222 U145 ( .A(n90), .B(B[6]), .C(n57), .D(n62), .Q(n56) );
  INV3 U146 ( .A(A[6]), .Q(n90) );
  CLKIN6 U147 ( .A(n64), .Q(n62) );
  NAND21 U148 ( .A(B[7]), .B(n181), .Q(n54) );
  INV0 U149 ( .A(A[7]), .Q(n181) );
  NAND22 U150 ( .A(B[8]), .B(net715532), .Q(n50) );
  INV3 U151 ( .A(A[8]), .Q(net715532) );
  NOR24 U152 ( .A(n93), .B(B[9]), .Q(n47) );
  NAND21 U153 ( .A(B[9]), .B(n93), .Q(n48) );
  INV3 U154 ( .A(A[9]), .Q(n93) );
  NOR23 U155 ( .A(n17), .B(n28), .Q(n15) );
  INV2 U156 ( .A(n184), .Q(n190) );
  INV6 U157 ( .A(n30), .Q(n184) );
  NOR22 U158 ( .A(n38), .B(n40), .Q(n36) );
  NOR24 U159 ( .A(n180), .B(B[11]), .Q(n38) );
  NOR21 U160 ( .A(n179), .B(B[10]), .Q(n40) );
  INV3 U161 ( .A(A[10]), .Q(n179) );
  NOR24 U162 ( .A(n31), .B(n185), .Q(n29) );
  OAI212 U163 ( .A(n32), .B(n35), .C(n33), .Q(n31) );
  NAND22 U164 ( .A(B[12]), .B(net715564), .Q(n35) );
  INV3 U165 ( .A(A[12]), .Q(net715564) );
  NOR24 U166 ( .A(n182), .B(B[13]), .Q(n32) );
  NAND21 U167 ( .A(B[13]), .B(n182), .Q(n33) );
  INV3 U168 ( .A(A[13]), .Q(n182) );
  NOR24 U169 ( .A(n184), .B(n183), .Q(n185) );
  OAI212 U170 ( .A(n38), .B(n41), .C(n39), .Q(n37) );
  NAND23 U171 ( .A(B[10]), .B(n179), .Q(n41) );
  NAND21 U172 ( .A(B[11]), .B(n180), .Q(n39) );
  INV3 U173 ( .A(A[11]), .Q(n180) );
  NOR23 U174 ( .A(n23), .B(n19), .Q(n18) );
  OAI212 U175 ( .A(n27), .B(n24), .C(n25), .Q(n23) );
  NAND22 U176 ( .A(B[14]), .B(net715472), .Q(n27) );
  INV3 U177 ( .A(A[14]), .Q(net715472) );
  NOR24 U178 ( .A(n178), .B(B[15]), .Q(n24) );
  NAND21 U179 ( .A(B[15]), .B(n178), .Q(n25) );
  INV3 U180 ( .A(A[15]), .Q(n178) );
  NAND24 U181 ( .A(n20), .B(n21), .Q(n19) );
  NOR24 U182 ( .A(n189), .B(n186), .Q(n188) );
  CLKIN6 U183 ( .A(n7), .Q(n189) );
  NOR24 U184 ( .A(n8), .B(n11), .Q(n7) );
  NAND24 U185 ( .A(n10), .B(n9), .Q(n8) );
  NOR22 U186 ( .A(B[24]), .B(B[25]), .Q(n10) );
  NOR23 U187 ( .A(B[26]), .B(B[27]), .Q(n9) );
  NAND24 U188 ( .A(n12), .B(n13), .Q(n11) );
  NOR22 U189 ( .A(B[23]), .B(B[22]), .Q(n12) );
  NOR23 U190 ( .A(B[21]), .B(B[20]), .Q(n13) );
  NOR23 U191 ( .A(B[30]), .B(n4), .Q(n3) );
  NAND24 U192 ( .A(n6), .B(n5), .Q(n4) );
  INV3 U193 ( .A(B[28]), .Q(n6) );
  INV3 U194 ( .A(B[29]), .Q(n5) );
  NOR24 U195 ( .A(n90), .B(B[6]), .Q(n59) );
  NOR22 U196 ( .A(n24), .B(n26), .Q(n22) );
  NOR22 U197 ( .A(net715472), .B(B[14]), .Q(n26) );
  NOR24 U198 ( .A(net715318), .B(B[3]), .Q(n76) );
  NOR24 U199 ( .A(net715564), .B(B[12]), .Q(n34) );
  CLKIN6 U200 ( .A(n76), .Q(n74) );
  NOR24 U201 ( .A(n34), .B(n32), .Q(n30) );
  NOR23 U202 ( .A(net715532), .B(B[8]), .Q(n49) );
endmodule


module sqroot_comb_NBITS32 ( arg, roundup, sqroot );
  input [31:0] arg;
  output [16:0] sqroot;
  input roundup;
  wire   res_31_, res_30_, res_29_, res_28_, res_27_, res_26_, res_25_,
         res_24_, res_23_, res_22_, res_21_, res_20_, res_19_, res_17_,
         res_16_, res_15_, res_14_, res_13_, res_12_, res_11_, res_10_, res_9_,
         res_8_, res_7_, res_6_, res_5_, res_4_, res_3_, res_2_, res_1_,
         res_0_, N1776, N1777, N1779, N1780, N1781, N1782, N1783, N1784, N1785,
         N1786, N1788, N1790, N1793, N1794, N1893, N1894, N1895, N1896, N1897,
         N1898, N1899, N1900, N1901, N1902, N1903, N1904, N1905, N1906, N1907,
         N1908, N1909, N1910, N1911, N1912, N1913, N1914, N1915, N1916, N1917,
         N1918, N1919, N1920, N1921, N1922, N1923, N1924, N1964, N1968, N1971,
         N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981, N1983,
         N1985, N1986, N1987, N2085, N2086, N2087, N2088, N2089, N2090, N2091,
         N2092, N2093, N2094, N2095, N2096, N2097, N2098, N2099, N2100, N2101,
         N2102, N2103, N2104, N2105, N2106, N2107, N2108, N2109, N2110, N2111,
         N2112, N2113, N2114, N2115, N2116, N2243, N2277, N2278, N2279, N2280,
         N2281, N2282, N2283, N2284, N2285, N2286, N2287, N2288, N2289, N2290,
         N2291, N2292, N2293, N2294, N2295, N2296, N2297, N2298, N2299, N2300,
         N2301, N2302, N2303, N2304, N2305, N2306, N2307, N2308, N2435, N2474,
         N2475, N2476, N2477, N2478, N2479, N2480, N2481, N2482, N2483, N2484,
         N2485, N2486, N2487, N2488, N2489, N2490, N2491, N2492, N2493, N2494,
         N2495, N2496, N2497, N2498, N2499, N2500, N2538, N2540, N2541, N2542,
         N2543, N2544, N2545, N2546, N2548, N2549, N2550, N2551, N2552, N2553,
         N2554, N2556, N2557, N2559, N2560, N2561, N2627, N2661, N2662, N2663,
         N2664, N2665, N2666, N2667, N2668, N2669, N2670, N2671, N2672, N2673,
         N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682, N2683,
         N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692, N2819,
         N2854, N2855, N2856, N2857, N2858, N2859, N2860, N2861, N2862, N2863,
         N2864, N2865, N2866, N2867, N2868, N2869, N2870, N2871, N2872, N2873,
         N2874, N2875, N2876, N2877, N2878, N2879, N2880, N2881, N2882, N2883,
         N2884, N2947, N2950, N2951, N2952, N2953, N2954, N2955, N2956, N2957,
         N2958, N2959, N2960, N2961, N2962, N2963, N2964, N2965, N2966,
         net640122, N2063, net660260, net660303, net660309, net675324,
         net702066, net703634, net703782, net703797, net710022, net711876,
         net711884, net711901, net711939, net711940, net712018, net712020,
         net712079, net712089, net712113, net712114, net712123, net712124,
         net712125, net712126, net712127, net712129, net712130, net712132,
         net712133, net712134, net712139, net712145, net712146, net712147,
         net712148, net712151, net712164, net712165, net712166, net712167,
         net712168, net712169, net712171, net712175, net712196, net712197,
         net712199, net712202, net712203, net712208, net712211, net712214,
         net712216, net712238, net712286, net712305, net712307, net712311,
         net712316, net712323, net712328, net712330, net712341, net712344,
         net712357, net712359, net712361, net712363, net712366, net712369,
         net712374, net712410, net712412, net712414, net712415, net712433,
         net712434, net712454, net712460, net712461, net712462, net712475,
         net712478, net712483, net712484, net712493, net712496, net712501,
         net712502, net712503, net712504, net712505, net712507, net712512,
         net712513, net712518, net712521, net712529, net712531, net712535,
         net712536, net712544, net712555, net712559, net712560, net712567,
         net712568, net712569, net712573, net712582, net712587, net712588,
         net712595, net712596, net712600, net712602, net712605, net712610,
         net712612, net712619, net712620, net712634, net712637, net712642,
         net712644, net712646, net712651, net712652, net712654, net712655,
         net712656, net712668, net712672, net712674, net712677, net712680,
         net712688, net712696, net712698, net712700, net712702, net712704,
         net712710, net712712, net712716, net712721, net712722, net712727,
         net712729, net712730, net712731, net712732, net712733, net712743,
         net712744, net712746, net712751, net712752, net712753, net712754,
         net712755, net712760, net712766, net712773, net712774, net712775,
         net712777, net712778, net712781, net712782, net712784, net712787,
         net712788, net712789, net712790, net712792, net712793, net712803,
         net712810, net712815, net712816, net712819, net712821, net712824,
         net712825, net712831, net712842, net712848, net712855, net712860,
         net712864, net712865, net712871, net712877, net712879, net712880,
         net712881, net712885, net712887, net712888, net712893, net712894,
         net712895, net712898, net712899, net712901, net712902, net712903,
         net712904, net712905, net712910, net712914, net712917, net712918,
         net712919, net712929, net712931, net712934, net712935, net712938,
         net712939, net712940, net712941, net712945, net712946, net712950,
         net712951, net712952, net712957, net712959, net712960, net712963,
         net712965, net712966, net712967, net712970, net712976, net712977,
         net712979, net712980, net712983, net712984, net712985, net712990,
         net712991, net712992, net712993, net712996, net712997, net713001,
         net713002, net713005, net713008, net713009, net713011, net713015,
         net713020, net713024, net713031, net713041, net713043, net713044,
         net713045, net713047, net713051, net713052, net713053, net713055,
         net713057, net713058, net713061, net713066, net713067, net713068,
         net713072, net713073, net713074, net713078, net713084, net713085,
         net713087, net713090, net713096, net713097, net713098, net713099,
         net713100, net713101, net713103, net713104, net713114, net713116,
         net713125, net713127, net713129, net713130, net713138, net713141,
         net713142, net713143, net713146, net713148, net713149, net713150,
         net713151, net713152, net713153, net713155, net713157, net713158,
         net713159, net713160, net713161, net713162, net713166, net713167,
         net713169, net713170, net713171, net713181, net713184, net713186,
         net713189, net713193, net713194, net713196, net713197, net713199,
         net713210, net713211, net715326, net715348, net715346, net715344,
         net715362, net715360, net715376, net715416, net715412, net715406,
         net715402, net715450, net715480, net715478, net715510, net715506,
         net715544, net715542, net715540, net715576, net715572, net715570,
         net715616, net715614, net715610, net715608, net715606, net715680,
         net715678, net715674, net715687, net715700, net715705, net715704,
         net715712, net715711, net715710, net715719, net715717, net715725,
         net715739, net715746, net715745, net715754, net715753, net715761,
         net715759, net715769, net715768, net715767, net715766, net715776,
         net715775, net715783, net715782, net715781, net715788, net715794,
         net715804, net715803, net715802, net715816, net715825, net715824,
         net716101, net716133, net716172, net716181, net716206, net716222,
         net716268, net716366, net716390, net716389, net716402, net716401,
         net716699, net717453, net717664, net717806, net717816, net717815,
         net717814, net717907, net718011, net718067, net718090, net718129,
         net718128, net718162, net718226, net718324, net718339, net718343,
         net718362, net718373, net718388, net718432, net718447, net718466,
         net718473, net718471, net718490, net718495, net718535, net718534,
         net718580, net718604, net718619, net718618, net718617, net718624,
         net719152, net719166, net719165, net719234, net719237, net719293,
         net719298, net719306, net719327, net719447, net719548, net719603,
         net719607, net719606, net719616, net719615, net719727, net719733,
         net719772, net719771, net719953, net719952, net719966, net719965,
         net719964, net720042, net720041, net720124, net720121, net720185,
         net720253, net720274, net720318, net720325, net720329, net720403,
         net720401, net720567, net720570, net720700, net720699, net720697,
         net720693, net720727, net720783, net720787, net720826, net720894,
         net720951, net720967, net720986, net721014, net721024, net721034,
         net721041, net721083, net721078, net721077, net721134, net721162,
         net721166, net721242, net721256, net721268, net721293, net721315,
         net721341, net721340, net721349, net721373, net721379, net721406,
         net721440, net721443, net721548, net721638, net721637, net721629,
         net721714, net721808, net721834, net722174, net722205, net722204,
         net722223, net722222, net722234, net722399, net722414, net722413,
         net722422, net722433, net722482, net722521, net722561, net722560,
         net722729, net722738, net722889, net722912, net723106, net723109,
         net723251, net723273, net723292, net723417, net723419, net723431,
         net723435, net723444, net723472, net723480, net723498, net723514,
         net723527, net723538, net723541, net723547, net723555, net723577,
         net723603, net723620, net723637, net723674, net723702, net723742,
         net723751, net723758, net723768, net723781, net723850, net723873,
         net723881, net723883, net723890, net723891, net723912, net723918,
         net723917, net723927, net723959, net723961, net723969, net724003,
         net724008, net724021, net724065, net724072, net724116, net724119,
         net724125, net724167, net724188, net724284, net724374, net724429,
         net724508, net724566, net724671, net724738, net724758, net724789,
         net724795, net724837, net724864, net724863, net724923, net724932,
         net725117, net725181, net725214, net725420, net725419, net725440,
         net725448, net725453, net725460, net725473, net725472, net725476,
         net725513, net725636, net725635, net725641, net725733, net725903,
         net725944, net726021, net726092, net726138, net726169, net726168,
         net726165, net726276, net726353, net715646, net715642, net712607,
         net706857, net715508, net712758, net712589, net725046, net713118,
         net713117, net713112, net713109, net712942, net712804, net725112,
         net713121, net713120, net713102, net713046, net726012, net721410,
         net721408, net712184, net712087, net712190, net712189, net712188,
         net712186, net712192, net712131, net716332, net716331, net711990,
         net711886, net715378, net715374, N2547, n2862, n2863, n2864, n2865,
         n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875,
         n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885,
         n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895,
         n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905,
         n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915,
         n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925,
         n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935,
         n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945,
         n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955,
         n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965,
         n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975,
         n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985,
         n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995,
         n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025,
         n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035,
         n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045,
         n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055,
         n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065,
         n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075,
         n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085,
         n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095,
         n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105,
         n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115,
         n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125,
         n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135,
         n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145,
         n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155,
         n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165,
         n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175,
         n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185,
         n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195,
         n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205,
         n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215,
         n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225,
         n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255,
         n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265,
         n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275,
         n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285,
         n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295,
         n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305,
         n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315,
         n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325,
         n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335,
         n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345,
         n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355,
         n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365,
         n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375,
         n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385,
         n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395,
         n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405,
         n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415,
         n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425,
         n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435,
         n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445,
         n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455,
         n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
         n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
         n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
         n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
         n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
         n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
         n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
         n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
         n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
         n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
         n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
         n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
         n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
         n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
         n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
         n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
         n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
         n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
         n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
         n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
         n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
         n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
         n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
         n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
         n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
         n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
         n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
         n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
         n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
         n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
         n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
         n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
         n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
         n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
         n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
         n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
         n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
         n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
         n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
         n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
         n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
         n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, SYNOPSYS_UNCONNECTED_1,
         SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3,
         SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5,
         SYNOPSYS_UNCONNECTED_6;

  sqroot_comb_NBITS32_DW01_sub_28 sub_0_root_sub_0_root_sub_44_I15 ( .A({n3502, 
        n3505, n3542, N2560, N2559, n3454, n3347, N2556, n3517, N2554, N2553, 
        n3540, N2551, N2550, N2549, n3555, net716366, N2546, N2545, N2544, 
        n3541, n3249, n3203, n3350, n3400, N2538, n3258, n4233, n4235, n3530, 
        n4234, n3232}), .B({n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, net715775, net715783, 
        net715825, net715803, net715606, net715788, net725733, net715794, 
        net716133, net726169, net715761, n3575, net715725, net719306, n4257, 
        n4256, n4257, n4257}), .CI(n4257), .DIFF({N2692, N2691, N2690, N2689, 
        N2688, N2687, N2686, N2685, N2684, N2683, N2682, N2681, N2680, N2679, 
        N2678, N2677, N2676, N2675, N2674, N2673, N2672, N2671, N2670, N2669, 
        N2668, N2667, N2666, N2665, N2664, N2663, N2662, N2661}) );
  sqroot_comb_NBITS32_DW01_inc_3 add_53 ( .A({n4257, net715775, net715781, 
        net725513, net715802, net715606, net715788, net725733, net715794, 
        net716133, net726169, net715761, n3576, net715725, net718226, 
        net723850, net720274}), .SUM({N2966, N2965, N2964, N2963, N2962, N2961, 
        N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, 
        N2950}) );
  sqroot_comb_NBITS32_DW01_sub_31 sub_0_root_sub_0_root_sub_44_I12 ( .A({N1987, 
        N1986, N1985, n3520, N1983, n3525, N1981, N1980, N1979, N1978, N1977, 
        N1976, N1975, N1974, N1973, net716268, N1971, n3230, net722738, N1968, 
        net722729, n3397, n3531, N1964, n3533, n3532, n3534, n3535, n3536, 
        n3538, n3537, n3539}), .B({n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, net715776, net715782, net715825, 
        net715804, net715606, net715788, net725733, net715794, net715816, 
        net724072, N2063, n4257, n4256, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257}), .CI(n4257), .DIFF({N2116, N2115, N2114, N2113, 
        N2112, N2111, N2110, N2109, N2108, N2107, N2106, N2105, N2104, N2103, 
        N2102, N2101, N2100, N2099, N2098, N2097, N2096, N2095, N2094, N2093, 
        N2092, N2091, N2090, N2089, N2088, N2087, N2086, N2085}) );
  sqroot_comb_NBITS32_DW01_sub_32 sub_0_root_sub_0_root_sub_44_I11 ( .A({n4226, 
        N1794, n3285, n3192, n3527, N1790, n3506, N1788, n3333, N1786, N1785, 
        N1784, N1783, N1782, N1781, N1780, N1779, n3529, N1777, N1776, 
        arg[11:0]}), .B({n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, net715775, net715782, net725513, net715802, 
        net715606, net715788, net724508, net715794, net715816, net715700, 
        n4257, n4256, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257}), .CI(n4257), .DIFF({N1924, N1923, N1922, N1921, N1920, 
        N1919, N1918, N1917, N1916, N1915, N1914, N1913, N1912, N1911, N1910, 
        N1909, N1908, N1907, N1906, N1905, N1904, N1903, N1902, N1901, N1900, 
        N1899, N1898, N1897, N1896, N1895, N1894, N1893}) );
  sqroot_comb_NBITS32_DW01_sub_39 sub_0_root_sub_0_root_sub_44_I13 ( .A({n3226, 
        n3228, n4255, n3524, n3339, n3523, n3514, n2926, n4254, n4253, n4252, 
        n3513, n3231, net660260, n4251, n3227, n3264, n4250, n3522, net725214, 
        n3327, n2925, n3239, n3528, n4292, n4293, n4294, n4295, n4296, n4297, 
        n4298, n4299}), .B({n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, net715776, net715782, net725513, 
        net715804, net715606, net715788, net725733, net715794, net716133, 
        net726169, net715761, n3575, n4257, n4256, n4257, n4257, n4257, n4257, 
        n4257, n4257}), .CI(n4257), .DIFF({N2308, N2307, N2306, N2305, N2304, 
        N2303, N2302, N2301, N2300, N2299, N2298, N2297, N2296, N2295, N2294, 
        N2293, N2292, N2291, N2290, N2289, N2288, N2287, N2286, N2285, N2284, 
        N2283, N2282, N2281, N2280, N2279, N2278, N2277}) );
  sqroot_comb_NBITS32_DW01_sub_43 sub_1_root_sub_44_I16 ( .A({n4258, n4216, 
        n4224, n4261, n4262, n4218, n4221, n4213, n4215, n4217, n4220, n4212, 
        n4214, n4222, n3277, n3552, n3439, n4275, net640122, n3548, n3550, 
        n4278, n4279, n3551, n3544, n4282, n3423, net703797, n3545, n4285, 
        n3546, n4232}), .B({n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, net715775, 
        net715781, net715824, net715802, net715606, net715788, net725733, 
        net715794, net715816, net726169, net715761, n3576, net715725, 
        net725641, net717664, n4257, n4257}), .CI(n4256), .DIFF({N2884, N2883, 
        N2882, N2881, N2880, N2879, N2878, N2877, N2876, N2875, N2874, N2873, 
        N2872, N2871, N2870, N2869, N2868, N2867, N2866, N2865, N2864, N2863, 
        N2862, N2861, N2860, N2859, N2858, N2857, N2856, N2855, N2854, 
        SYNOPSYS_UNCONNECTED_1}) );
  sqroot_comb_NBITS32_DW_cmp_45 lte_43_I13 ( .A({n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, net715775, 
        net715783, net715825, net715802, net715606, net715788, net725733, 
        net715794, net716133, net726169, net715761, n3576, n4257, n4256, n4257, 
        n4257, n4257, n4257, n4257, n4257}), .B({n3226, n3228, n4255, n3524, 
        n3339, n3523, n3514, n2926, n4254, n4253, n4252, n3513, n3231, 
        net660260, n4251, n3227, n3264, n4250, n3522, net725214, n3305, n2925, 
        n3239, n3528, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299}), 
        .TC(n4257), .GE_LT(n4257), .GE_GT_EQ(n4257), .GE_LT_GT_LE(N2243) );
  sqroot_comb_NBITS32_DW_cmp_47 lte_43_I15 ( .A({n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        net715775, net715783, net725513, net715803, net715606, net715788, 
        net725733, net715794, net716133, net726169, net715761, n3576, 
        net715725, net718129, n4257, n4256, n4257, n4257}), .B({n3502, n3505, 
        n3542, N2560, N2559, n3454, n3347, N2556, n3517, N2554, N2553, n3540, 
        N2551, N2550, N2549, N2548, net716366, N2546, N2545, N2544, n3541, 
        n3249, n3203, N2540, n3400, n3554, n3258, n4233, n4235, n3530, n4234, 
        n3232}), .TC(n4257), .GE_LT(n4257), .GE_GT_EQ(n4257), .GE_LT_GT_LE(
        N2627) );
  sqroot_comb_NBITS32_DW_cmp_49 lte_43_I14 ( .A({n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        net715776, net715781, net715824, net715804, net715606, net715788, 
        net715704, net715794, net716133, net726169, net715761, n3576, 
        net723969, n4257, n4256, n4257, n4257, n4257, n4257}), .B({n3519, 
        n3229, n4249, n3262, n4248, n3518, n4247, n4246, n3521, n3440, n4245, 
        n3261, n3298, n4230, n4227, n4228, net660303, n4244, n4243, net660309, 
        n4242, n4241, n4240, n4239, n3516, n4238, n4237, n4236, n4235, n3530, 
        n4234, n3232}), .TC(n4257), .GE_LT(n4257), .GE_GT_EQ(n4257), 
        .GE_LT_GT_LE(N2435) );
  sqroot_comb_NBITS32_DW_cmp_50 lte_43_I16 ( .A({n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, net715775, net715782, net715825, net715803, net715606, 
        net715788, net725733, net715794, net716133, net726169, net715761, 
        n3575, net715725, net718226, net715739, n4257, n4256}), .B({n4258, 
        n4259, n4260, n3247, n4231, n4263, n4264, n4265, n4266, n4267, n4268, 
        n4269, n4270, n4271, n4272, n3552, n4274, n4275, net640122, n3548, 
        n3550, n4223, n4211, n3551, n3544, n4282, n4283, net703797, n3545, 
        n4219, n3437, n4287}), .TC(n4257), .GE_LT(n4257), .GE_GT_EQ(n4257), 
        .GE_LT_GT_LE(N2819) );
  sqroot_comb_NBITS32_DW01_sub_69 sub_0_root_sub_0_root_sub_44_I14 ( .A({n3519, 
        n3229, n4249, n3262, n4248, n3518, n4247, n4246, n3521, n3440, n4245, 
        n3261, n3298, n4288, n4289, n4290, net660303, n4244, n4243, net660309, 
        n4291, n3418, n4240, n4239, n3516, n4238, n4237, n4236, n4235, n3530, 
        n4234, n3232}), .B({n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, net715776, net715783, 
        net725513, net715804, net715606, net715788, net725733, net715794, 
        net716133, net726169, net715761, n3575, net715719, n4257, n4256, n4257, 
        n4257, n4257, n4257}), .CI(n4257), .DIFF({N2500, N2499, N2498, N2497, 
        N2496, N2495, N2494, N2493, N2492, N2491, N2490, N2489, N2488, N2487, 
        N2486, N2485, N2484, N2483, N2482, N2481, N2480, N2479, N2478, N2477, 
        N2476, N2475, N2474, SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, 
        SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6}) );
  sqroot_comb_NBITS32_DW_cmp_48 lt_gt_52 ( .A({n4257, n4257, n4257, n4257, 
        n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, n4257, 
        n4257, n4257, net715775, net715781, net725513, net715803, net715606, 
        net715788, net725733, net715794, net716133, net726169, net715761, 
        n3575, net715725, net718226, net724671, net715754}), .B({res_31_, 
        res_30_, res_29_, res_28_, res_27_, res_26_, res_25_, res_24_, res_23_, 
        res_22_, res_21_, res_20_, res_19_, n4229, res_17_, res_16_, res_15_, 
        res_14_, res_13_, res_12_, res_11_, res_10_, res_9_, res_8_, res_7_, 
        res_6_, res_5_, res_4_, res_3_, res_2_, res_1_, res_0_}), .TC(n4257), 
        .GE_LT(n4256), .GE_GT_EQ(n4257), .GE_LT_GT_LE(N2947) );
  NAND24 U2842 ( .A(net712568), .B(net723912), .Q(net712366) );
  NAND26 U2843 ( .A(n3774), .B(n3252), .Q(net712568) );
  CLKIN8 U2844 ( .A(net717664), .Q(net721041) );
  CLKIN2 U2845 ( .A(n4275), .Q(n4190) );
  BUF2 U2846 ( .A(n3258), .Q(n2862) );
  BUF2 U2847 ( .A(n3440), .Q(n2863) );
  INV15 U2848 ( .A(net715344), .Q(net719327) );
  INV12 U2849 ( .A(net723620), .Q(net718324) );
  NAND21 U2850 ( .A(N2490), .B(net723620), .Q(n4083) );
  INV4 U2851 ( .A(net719293), .Q(net719298) );
  NAND23 U2852 ( .A(n3801), .B(net715616), .Q(net712704) );
  XOR22 U2853 ( .A(n2929), .B(n3156), .Q(net723431) );
  NAND34 U2854 ( .A(n3836), .B(n3835), .C(n3929), .Q(n3476) );
  NAND24 U2855 ( .A(n3796), .B(n3186), .Q(n3835) );
  INV6 U2856 ( .A(net712462), .Q(net712369) );
  CLKIN12 U2857 ( .A(net715646), .Q(net726021) );
  INV8 U2858 ( .A(net712535), .Q(net723273) );
  NOR23 U2859 ( .A(n2905), .B(n2906), .Q(n2907) );
  OAI210 U2860 ( .A(arg[13]), .B(net723637), .C(net716172), .Q(n3922) );
  NAND23 U2861 ( .A(n2914), .B(n3997), .Q(n3909) );
  OAI211 U2862 ( .A(n3877), .B(n3876), .C(n3875), .Q(n3994) );
  NAND22 U2863 ( .A(n3204), .B(net712475), .Q(n3206) );
  NAND21 U2864 ( .A(n3540), .B(net719447), .Q(n4147) );
  NAND21 U2865 ( .A(N2550), .B(net719447), .Q(n4151) );
  NAND22 U2866 ( .A(n3325), .B(net719447), .Q(n4155) );
  NAND22 U2867 ( .A(n4138), .B(n4137), .Q(n4221) );
  AOI221 U2868 ( .A(n4132), .B(n4131), .C(net722560), .D(n4131), .Q(n3247) );
  BUF15 U2869 ( .A(net712559), .Q(net723912) );
  CLKIN6 U2870 ( .A(net712559), .Q(net712555) );
  INV2 U2871 ( .A(n3427), .Q(n3463) );
  NAND24 U2872 ( .A(net720041), .B(n3213), .Q(n3214) );
  CLKIN6 U2873 ( .A(n3696), .Q(n3480) );
  INV12 U2874 ( .A(net723768), .Q(net712607) );
  BUF12 U2875 ( .A(n3526), .Q(n3506) );
  INV2 U2876 ( .A(n3861), .Q(n2864) );
  NAND24 U2877 ( .A(net712521), .B(n3368), .Q(n3758) );
  OAI212 U2878 ( .A(net712139), .B(net716181), .C(n3832), .Q(n2865) );
  OAI211 U2879 ( .A(net712139), .B(net716181), .C(n3832), .Q(n3928) );
  NAND24 U2880 ( .A(n3197), .B(n3198), .Q(n3832) );
  AOI2111 U2881 ( .A(net721714), .B(net715816), .C(n3962), .D(n3961), .Q(n3966) );
  INV3 U2882 ( .A(n3920), .Q(n3962) );
  BUF2 U2883 ( .A(N1968), .Q(n2866) );
  INV8 U2884 ( .A(net712113), .Q(N1968) );
  NAND22 U2885 ( .A(net712199), .B(N1783), .Q(n3191) );
  BUF12 U2886 ( .A(net718129), .Q(n2867) );
  INV2 U2887 ( .A(net718162), .Q(net725440) );
  NAND23 U2888 ( .A(net725440), .B(n3217), .Q(n3218) );
  NAND22 U2889 ( .A(net725440), .B(n3300), .Q(n3483) );
  NAND26 U2890 ( .A(n3483), .B(n4110), .Q(n4275) );
  INV6 U2891 ( .A(net712203), .Q(N1973) );
  INV3 U2892 ( .A(n4002), .Q(n3990) );
  NAND26 U2893 ( .A(n2888), .B(n4002), .Q(n3915) );
  INV10 U2894 ( .A(n3973), .Q(N1783) );
  CLKIN6 U2895 ( .A(net712171), .Q(n2980) );
  NAND23 U2896 ( .A(net712214), .B(net715608), .Q(n3976) );
  NAND22 U2897 ( .A(net719298), .B(n4290), .Q(n3329) );
  INV3 U2898 ( .A(n2869), .Q(n3122) );
  BUF6 U2899 ( .A(net712803), .Q(net715704) );
  INV12 U2900 ( .A(net712567), .Q(net712634) );
  CLKIN15 U2901 ( .A(net712357), .Q(net712363) );
  NAND26 U2902 ( .A(n3487), .B(n3637), .Q(n3639) );
  NAND23 U2903 ( .A(n3650), .B(net712871), .Q(n3211) );
  INV4 U2904 ( .A(n3660), .Q(n3362) );
  CLKIN6 U2905 ( .A(net715705), .Q(n2871) );
  INV8 U2906 ( .A(net715704), .Q(net712139) );
  INV12 U2907 ( .A(n3246), .Q(n3661) );
  NAND28 U2908 ( .A(net718373), .B(net712976), .Q(n3490) );
  CLKIN10 U2909 ( .A(net712819), .Q(net724008) );
  NAND26 U2910 ( .A(net721166), .B(net715767), .Q(n2868) );
  NAND24 U2911 ( .A(net721166), .B(net715767), .Q(net712819) );
  NAND23 U2912 ( .A(n3735), .B(net723912), .Q(n3745) );
  NAND22 U2913 ( .A(net722738), .B(net715544), .Q(n4021) );
  NAND22 U2914 ( .A(n3092), .B(n3134), .Q(n2942) );
  OAI211 U2915 ( .A(n3935), .B(n3415), .C(n3930), .Q(n3844) );
  NAND26 U2916 ( .A(net718473), .B(net712018), .Q(N2545) );
  INV8 U2917 ( .A(net712941), .Q(net712957) );
  CLKIN2 U2918 ( .A(net713143), .Q(net713155) );
  INV8 U2919 ( .A(net712816), .Q(net719152) );
  NAND24 U2920 ( .A(net712860), .B(net723435), .Q(n2869) );
  NAND28 U2921 ( .A(n3489), .B(n3490), .Q(net712860) );
  CLKIN3 U2922 ( .A(n3789), .Q(n3204) );
  CLKIN3 U2923 ( .A(n3792), .Q(n3196) );
  BUF2 U2924 ( .A(net712359), .Q(n2934) );
  NAND23 U2925 ( .A(net712652), .B(net721373), .Q(n3776) );
  INV6 U2926 ( .A(net712743), .Q(net712754) );
  AOI222 U2927 ( .A(arg[17]), .B(net712787), .C(n2939), .D(net712139), .Q(
        net712784) );
  IMUX24 U2928 ( .A(net712959), .B(net712960), .S(n2870), .Q(n3631) );
  XNR21 U2929 ( .A(n3275), .B(arg[23]), .Q(n2870) );
  CLKIN6 U2930 ( .A(n2871), .Q(n2872) );
  BUF6 U2931 ( .A(net712792), .Q(net715705) );
  BUF6 U2932 ( .A(net715506), .Q(n2873) );
  NAND26 U2933 ( .A(n3631), .B(n3496), .Q(net712848) );
  NAND26 U2934 ( .A(n2957), .B(n2958), .Q(net712696) );
  NAND28 U2935 ( .A(n3646), .B(net715608), .Q(n3657) );
  NAND26 U2936 ( .A(net712792), .B(n3109), .Q(n3108) );
  NAND26 U2937 ( .A(n3649), .B(net712803), .Q(n3650) );
  NAND23 U2938 ( .A(n3927), .B(net721637), .Q(n3335) );
  NAND26 U2939 ( .A(n3219), .B(n3623), .Q(n3444) );
  CLKIN6 U2940 ( .A(n3365), .Q(n3643) );
  INV6 U2941 ( .A(net712980), .Q(net712979) );
  NAND24 U2942 ( .A(n3659), .B(net712792), .Q(n3660) );
  NAND23 U2943 ( .A(net712286), .B(n3926), .Q(n3927) );
  BUF2 U2944 ( .A(n3724), .Q(n2874) );
  INV0 U2945 ( .A(net723751), .Q(net722174) );
  INV3 U2946 ( .A(net725944), .Q(n2978) );
  CLKBU15 U2947 ( .A(n3889), .Q(n2895) );
  INV3 U2948 ( .A(n3661), .Q(n3442) );
  NAND24 U2949 ( .A(n3996), .B(n3293), .Q(N1794) );
  INV6 U2950 ( .A(N1923), .Q(n4024) );
  INV0 U2951 ( .A(n4018), .Q(n2875) );
  CLKIN3 U2952 ( .A(net719771), .Q(net719772) );
  INV3 U2953 ( .A(n3397), .Q(n4018) );
  NAND26 U2954 ( .A(n2921), .B(net712192), .Q(net712131) );
  INV10 U2955 ( .A(n3958), .Q(n4014) );
  BUF2 U2956 ( .A(net716699), .Q(n2876) );
  CLKIN8 U2957 ( .A(net721014), .Q(net716699) );
  CLKIN12 U2958 ( .A(net723109), .Q(net712778) );
  NAND28 U2959 ( .A(n3326), .B(net712781), .Q(net723109) );
  NAND28 U2960 ( .A(n3488), .B(n3645), .Q(n3279) );
  CLKIN15 U2961 ( .A(net712589), .Q(net712758) );
  INV1 U2962 ( .A(net712729), .Q(net712751) );
  NAND22 U2963 ( .A(net716389), .B(net715781), .Q(n3392) );
  INV12 U2964 ( .A(n3943), .Q(n3970) );
  INV3 U2965 ( .A(n3344), .Q(n4020) );
  INV10 U2966 ( .A(n3722), .Q(n3414) );
  NAND21 U2967 ( .A(n2869), .B(n3467), .Q(n2877) );
  NAND22 U2968 ( .A(n2878), .B(n2879), .Q(n2880) );
  NAND23 U2969 ( .A(n2880), .B(n4198), .Q(res_9_) );
  INV2 U2970 ( .A(net715754), .Q(n2878) );
  INV3 U2971 ( .A(n4199), .Q(n2879) );
  INV2 U2972 ( .A(n4211), .Q(n4199) );
  NAND24 U2973 ( .A(net713068), .B(net713067), .Q(n3432) );
  NAND26 U2974 ( .A(n2993), .B(net713087), .Q(n2992) );
  NAND28 U2975 ( .A(net713066), .B(net715572), .Q(net712935) );
  INV6 U2976 ( .A(net724003), .Q(net721379) );
  INV6 U2977 ( .A(net712825), .Q(net720697) );
  NAND26 U2978 ( .A(n3447), .B(n3448), .Q(net712700) );
  CLKIN12 U2979 ( .A(n3296), .Q(n3219) );
  NAND26 U2980 ( .A(net720727), .B(n3411), .Q(n3413) );
  CLKIN4 U2981 ( .A(net712848), .Q(net712918) );
  NAND21 U2982 ( .A(net724738), .B(net712902), .Q(n3046) );
  NAND22 U2983 ( .A(net724738), .B(net712997), .Q(n3052) );
  NAND26 U2984 ( .A(net713072), .B(net713074), .Q(net703782) );
  INV4 U2985 ( .A(net713058), .Q(n3070) );
  CLKIN8 U2986 ( .A(n3063), .Q(n3087) );
  NAND22 U2987 ( .A(arg[21]), .B(net712979), .Q(n2882) );
  NAND22 U2988 ( .A(net712980), .B(n2881), .Q(n2883) );
  NAND24 U2989 ( .A(n2882), .B(n2883), .Q(n3646) );
  INV3 U2990 ( .A(arg[21]), .Q(n2881) );
  INV8 U2991 ( .A(net722413), .Q(net722414) );
  NAND26 U2992 ( .A(n3497), .B(n3618), .Q(n3619) );
  NAND28 U2993 ( .A(n3412), .B(n3413), .Q(n3618) );
  NAND32 U2994 ( .A(net713151), .B(n2896), .C(net713150), .Q(net713193) );
  INV10 U2995 ( .A(net713158), .Q(net713142) );
  NAND21 U2996 ( .A(N1918), .B(net715402), .Q(n4046) );
  BUF2 U2997 ( .A(net715402), .Q(net715759) );
  OAI212 U2998 ( .A(arg[11]), .B(net716101), .C(net715406), .Q(n4017) );
  INV12 U2999 ( .A(net715406), .Q(net715402) );
  CLKIN10 U3000 ( .A(n2974), .Q(net660309) );
  CLKIN15 U3001 ( .A(net716206), .Q(net725944) );
  INV6 U3002 ( .A(n3006), .Q(n2990) );
  INV2 U3003 ( .A(N1913), .Q(n2975) );
  NAND24 U3004 ( .A(n2886), .B(n2887), .Q(n2888) );
  INV6 U3005 ( .A(n4277), .Q(n3549) );
  INV12 U3006 ( .A(net723273), .Q(net723637) );
  NAND24 U3007 ( .A(n3611), .B(net715572), .Q(net713011) );
  INV6 U3008 ( .A(n3599), .Q(n3600) );
  NAND26 U3009 ( .A(n3724), .B(n3666), .Q(net712887) );
  NAND34 U3010 ( .A(net712130), .B(n4042), .C(net712129), .Q(net712127) );
  IMUX24 U3011 ( .A(n3328), .B(net723106), .S(n3578), .Q(n3327) );
  INV3 U3012 ( .A(net712199), .Q(net725903) );
  NAND34 U3013 ( .A(n2985), .B(net721408), .C(n2986), .Q(net721410) );
  MUX26 U3014 ( .A(net722738), .B(N2098), .S(n3575), .Q(n3522) );
  INV3 U3015 ( .A(net718011), .Q(net718067) );
  BUF6 U3016 ( .A(net718011), .Q(net723969) );
  INV6 U3017 ( .A(net712134), .Q(net712129) );
  INV4 U3018 ( .A(net722729), .Q(net726168) );
  NAND26 U3019 ( .A(n3763), .B(n3292), .Q(net712588) );
  INV0 U3020 ( .A(net726168), .Q(n2884) );
  NAND24 U3021 ( .A(n3209), .B(n3787), .Q(n3788) );
  CLKBU4 U3022 ( .A(net713116), .Q(n2897) );
  CLKIN6 U3023 ( .A(n3695), .Q(n3317) );
  INV6 U3024 ( .A(net712496), .Q(net712493) );
  BUF2 U3025 ( .A(n3140), .Q(net720318) );
  NAND34 U3026 ( .A(net712126), .B(net712125), .C(net712127), .Q(n2885) );
  INV6 U3027 ( .A(n3029), .Q(net712910) );
  NAND33 U3028 ( .A(net712126), .B(net712125), .C(net712127), .Q(net712124) );
  INV10 U3029 ( .A(net718534), .Q(net718535) );
  CLKIN4 U3030 ( .A(n3856), .Q(n3830) );
  CLKIN10 U3031 ( .A(net712484), .Q(net712535) );
  NAND26 U3032 ( .A(n3754), .B(net726021), .Q(n3755) );
  INV4 U3033 ( .A(n3575), .Q(n4054) );
  NAND28 U3034 ( .A(n3334), .B(net722912), .Q(n3336) );
  CLKIN6 U3035 ( .A(n3927), .Q(n3334) );
  CLKIN4 U3036 ( .A(n3944), .Q(n2886) );
  INV3 U3037 ( .A(net715769), .Q(n2887) );
  INV8 U3038 ( .A(n3092), .Q(n2941) );
  INV1 U3039 ( .A(net712361), .Q(net712344) );
  NAND22 U3040 ( .A(n3887), .B(net722889), .Q(n3865) );
  INV0 U3041 ( .A(net712544), .Q(n2889) );
  INV12 U3042 ( .A(net723577), .Q(net724374) );
  INV15 U3043 ( .A(net712286), .Q(net716172) );
  INV4 U3044 ( .A(net712501), .Q(n3170) );
  CLKIN3 U3045 ( .A(n3156), .Q(n2928) );
  NAND24 U3046 ( .A(n2928), .B(n2929), .Q(n2931) );
  NAND23 U3047 ( .A(n2959), .B(net719966), .Q(n3343) );
  NOR32 U3048 ( .A(n3460), .B(n3709), .C(net712716), .Q(n2890) );
  NAND26 U3049 ( .A(n3757), .B(net715678), .Q(n3748) );
  CLKIN10 U3050 ( .A(n3762), .Q(n3757) );
  NAND21 U3051 ( .A(N1920), .B(net715759), .Q(n4045) );
  NAND24 U3052 ( .A(n3866), .B(net715769), .Q(net712359) );
  INV4 U3053 ( .A(n3866), .Q(n2905) );
  INV12 U3054 ( .A(net712208), .Q(net716206) );
  INV12 U3055 ( .A(N2063), .Q(net712199) );
  IMUX20 U3056 ( .A(n2909), .B(n2891), .S(net711876), .Q(sqroot[11]) );
  INV15 U3057 ( .A(N2961), .Q(n2891) );
  INV0 U3058 ( .A(net703797), .Q(n2969) );
  NAND28 U3059 ( .A(n3834), .B(n3477), .Q(n3886) );
  NAND21 U3060 ( .A(n3314), .B(net723273), .Q(n3857) );
  CLKIN12 U3061 ( .A(net712361), .Q(n2892) );
  NAND24 U3062 ( .A(n3770), .B(n3216), .Q(net712569) );
  CLKIN6 U3063 ( .A(net715378), .Q(net715374) );
  CLKIN12 U3064 ( .A(net715378), .Q(net715376) );
  BUF2 U3065 ( .A(n3545), .Q(n2893) );
  NAND22 U3066 ( .A(N2483), .B(net723620), .Q(n4101) );
  NAND24 U3067 ( .A(n4101), .B(n4102), .Q(N2546) );
  BUF2 U3068 ( .A(n2875), .Q(n2894) );
  CLKIN3 U3069 ( .A(net713052), .Q(net713051) );
  NAND26 U3070 ( .A(n3082), .B(n3081), .Q(n3083) );
  INV6 U3071 ( .A(n3075), .Q(n3082) );
  NAND24 U3072 ( .A(n3075), .B(net713043), .Q(n3084) );
  NOR22 U3073 ( .A(net725944), .B(n3527), .Q(n4031) );
  NAND23 U3074 ( .A(N1916), .B(net725944), .Q(n4015) );
  NAND24 U3075 ( .A(n3619), .B(n3443), .Q(n3445) );
  OAI2112 U3076 ( .A(arg[26]), .B(n3017), .C(n3590), .D(arg[27]), .Q(n2896) );
  INV6 U3077 ( .A(net713031), .Q(net713116) );
  BUF2 U3078 ( .A(n3230), .Q(n2898) );
  BUF2 U3079 ( .A(n3227), .Q(n2899) );
  CLKIN6 U3080 ( .A(net718324), .Q(n2900) );
  CLKIN3 U3081 ( .A(n3987), .Q(n3571) );
  NAND22 U3082 ( .A(net712567), .B(net712357), .Q(net712560) );
  INV8 U3083 ( .A(net712704), .Q(net712596) );
  BUF12 U3084 ( .A(n3916), .Q(n3333) );
  CLKIN12 U3085 ( .A(net712605), .Q(net712619) );
  XNR21 U3086 ( .A(net715678), .B(net712781), .Q(n3707) );
  INV8 U3087 ( .A(n3080), .Q(net713072) );
  XNR22 U3088 ( .A(n3605), .B(net723480), .Q(n3606) );
  INV4 U3089 ( .A(n3899), .Q(n3902) );
  NAND22 U3090 ( .A(net725635), .B(net712366), .Q(n3899) );
  INV1 U3091 ( .A(n4005), .Q(n3390) );
  CLKIN12 U3092 ( .A(net712569), .Q(net712216) );
  CLKIN6 U3093 ( .A(n4072), .Q(n4064) );
  CLKIN6 U3094 ( .A(net713085), .Q(net713194) );
  NAND24 U3095 ( .A(net713129), .B(n3024), .Q(net713085) );
  NAND28 U3096 ( .A(net718339), .B(net712460), .Q(n2901) );
  NAND26 U3097 ( .A(net718339), .B(net712460), .Q(n3141) );
  NOR24 U3098 ( .A(n2907), .B(net712461), .Q(net712460) );
  OAI311 U3099 ( .A(n3603), .B(net713090), .C(net713143), .D(n3602), .Q(n3610)
         );
  NAND24 U3100 ( .A(n3220), .B(n3221), .Q(net712992) );
  NAND24 U3101 ( .A(net712934), .B(n3633), .Q(n3634) );
  INV4 U3102 ( .A(n3679), .Q(n3213) );
  INV6 U3103 ( .A(net712602), .Q(net712587) );
  NAND23 U3104 ( .A(n4012), .B(net724508), .Q(n3967) );
  BUF2 U3105 ( .A(n2926), .Q(n2902) );
  IMUX22 U3106 ( .A(N2102), .B(N1973), .S(net712079), .Q(n4057) );
  CLKIN0 U3107 ( .A(n2893), .Q(n4206) );
  NAND33 U3108 ( .A(n3314), .B(net723273), .C(n3315), .Q(n3316) );
  INV0 U3109 ( .A(n4251), .Q(n2903) );
  INV8 U3110 ( .A(n4057), .Q(n4251) );
  CLKIN8 U3111 ( .A(n2987), .Q(net660260) );
  NAND24 U3112 ( .A(net720042), .B(net720041), .Q(n3431) );
  INV3 U3113 ( .A(net723527), .Q(n3004) );
  INV10 U3114 ( .A(n3620), .Q(n3623) );
  INV15 U3115 ( .A(net712996), .Q(net718343) );
  NAND28 U3116 ( .A(n3647), .B(net715572), .Q(n3656) );
  CLKBU12 U3117 ( .A(n2873), .Q(net715788) );
  INV12 U3118 ( .A(net712919), .Q(net712831) );
  NAND28 U3119 ( .A(net712804), .B(net715768), .Q(net712919) );
  INV3 U3120 ( .A(net712721), .Q(net724789) );
  INV3 U3121 ( .A(net712722), .Q(net712721) );
  CLKIN6 U3122 ( .A(net712730), .Q(net723702) );
  NAND28 U3123 ( .A(n3815), .B(net715608), .Q(net724932) );
  NAND24 U3124 ( .A(net724932), .B(net712501), .Q(net712582) );
  NAND24 U3125 ( .A(net712710), .B(n2872), .Q(net712513) );
  INV1 U3126 ( .A(net723637), .Q(net716133) );
  INV10 U3127 ( .A(n3863), .Q(n3885) );
  NAND28 U3128 ( .A(n3472), .B(n3837), .Q(n3863) );
  CLKBU8 U3129 ( .A(net712199), .Q(net715406) );
  INV6 U3130 ( .A(net716268), .Q(net712196) );
  CLKIN12 U3131 ( .A(net712184), .Q(net726012) );
  INV15 U3132 ( .A(net719293), .Q(net722422) );
  NAND22 U3133 ( .A(n3902), .B(net712357), .Q(n3903) );
  BUF2 U3134 ( .A(n3722), .Q(n2904) );
  XNR20 U3135 ( .A(net721134), .B(n3736), .Q(n3779) );
  NAND24 U3136 ( .A(n4006), .B(n4005), .Q(n4007) );
  INV3 U3137 ( .A(n3282), .Q(n4006) );
  OAI211 U3138 ( .A(net720567), .B(n3569), .C(n3910), .Q(n3282) );
  NAND28 U3139 ( .A(net712573), .B(net715450), .Q(net712567) );
  NAND21 U3140 ( .A(n2868), .B(net712688), .Q(n3716) );
  XNR22 U3141 ( .A(net724566), .B(net712531), .Q(n3818) );
  CLKIN6 U3142 ( .A(net712374), .Q(net722889) );
  INV6 U3143 ( .A(net712410), .Q(net712374) );
  NAND23 U3144 ( .A(net702066), .B(net712702), .Q(n3696) );
  CLKIN4 U3145 ( .A(n3774), .Q(n3478) );
  CLKIN12 U3146 ( .A(n3688), .Q(n3326) );
  INV0 U3147 ( .A(net715768), .Q(n2906) );
  INV15 U3148 ( .A(net715766), .Q(net715768) );
  NAND24 U3149 ( .A(n4027), .B(n4026), .Q(n4028) );
  NAND21 U3150 ( .A(n3789), .B(net723891), .Q(n3205) );
  NAND28 U3151 ( .A(n2960), .B(net715616), .Q(net712855) );
  NAND26 U3152 ( .A(n3734), .B(net715540), .Q(net712656) );
  NAND22 U3153 ( .A(n3947), .B(n2909), .Q(n2910) );
  NAND26 U3154 ( .A(n2908), .B(net715606), .Q(n2911) );
  NAND24 U3155 ( .A(n2910), .B(n2911), .Q(n3948) );
  CLKIN6 U3156 ( .A(n3947), .Q(n2908) );
  CLKIN3 U3157 ( .A(net715606), .Q(n2909) );
  INV4 U3158 ( .A(n4010), .Q(N1788) );
  BUF2 U3159 ( .A(n3234), .Q(n2912) );
  INV0 U3160 ( .A(n3271), .Q(n2913) );
  INV1 U3161 ( .A(n3461), .Q(n3271) );
  CLKIN4 U3162 ( .A(n3821), .Q(n3461) );
  BUF4 U3163 ( .A(n3137), .Q(n2914) );
  INV6 U3164 ( .A(n3887), .Q(n2915) );
  INV2 U3165 ( .A(n3887), .Q(n3883) );
  INV10 U3166 ( .A(n3568), .Q(n3569) );
  CLKIN15 U3167 ( .A(n3663), .Q(n3687) );
  NAND43 U3168 ( .A(net724374), .B(net712595), .C(n3747), .D(n3269), .Q(n3268)
         );
  CLKIN4 U3169 ( .A(n3765), .Q(n3269) );
  INV12 U3170 ( .A(net712568), .Q(net720042) );
  CLKBU15 U3171 ( .A(n3886), .Q(n3236) );
  NAND23 U3172 ( .A(n3354), .B(net712504), .Q(n3797) );
  NAND22 U3173 ( .A(net722399), .B(net723890), .Q(n3354) );
  NAND23 U3174 ( .A(n3953), .B(n3952), .Q(n3954) );
  NAND22 U3175 ( .A(arg[12]), .B(net716172), .Q(n2918) );
  NAND24 U3176 ( .A(n2916), .B(n2917), .Q(n2919) );
  NAND28 U3177 ( .A(n2918), .B(n2919), .Q(N1776) );
  INV3 U3178 ( .A(arg[12]), .Q(n2916) );
  CLKIN3 U3179 ( .A(net716172), .Q(n2917) );
  NAND26 U3180 ( .A(net712196), .B(n2920), .Q(n2921) );
  INV0 U3181 ( .A(net715616), .Q(n2920) );
  NOR24 U3182 ( .A(net712131), .B(net712132), .Q(net712130) );
  NAND23 U3183 ( .A(n3214), .B(n3215), .Q(n3680) );
  INV3 U3184 ( .A(n3634), .Q(n3402) );
  INV2 U3185 ( .A(n3069), .Q(net724065) );
  CLKIN10 U3186 ( .A(n4100), .Q(n4233) );
  NAND23 U3187 ( .A(n3702), .B(net715572), .Q(net712722) );
  NAND22 U3188 ( .A(net718162), .B(N2667), .Q(n4119) );
  CLKIN6 U3189 ( .A(n3785), .Q(n3866) );
  INV6 U3190 ( .A(n2944), .Q(n2945) );
  INV6 U3191 ( .A(n3281), .Q(n3651) );
  CLKIN6 U3192 ( .A(n3788), .Q(n3810) );
  AOI2112 U3193 ( .A(n3772), .B(net723912), .C(net712560), .D(n2935), .Q(n3773) );
  NAND24 U3194 ( .A(arg[19]), .B(n3446), .Q(n3448) );
  NAND22 U3195 ( .A(net720697), .B(n3672), .Q(n2922) );
  NAND31 U3196 ( .A(n3682), .B(net723603), .C(n2923), .Q(net724003) );
  INV6 U3197 ( .A(n2922), .Q(n2923) );
  CLKIN4 U3198 ( .A(net721256), .Q(net723603) );
  CLKIN4 U3199 ( .A(net712483), .Q(net723918) );
  NAND24 U3200 ( .A(n3149), .B(net712238), .Q(n3147) );
  CLKIN10 U3201 ( .A(net712696), .Q(net712573) );
  NAND26 U3202 ( .A(net715642), .B(n3157), .Q(n3156) );
  INV1 U3203 ( .A(net717907), .Q(net718471) );
  NAND24 U3204 ( .A(N2477), .B(net717907), .Q(n3349) );
  INV6 U3205 ( .A(n4091), .Q(n3553) );
  NAND24 U3206 ( .A(n2951), .B(n2936), .Q(n2937) );
  NOR24 U3207 ( .A(net721834), .B(n3727), .Q(n3465) );
  CLKIN12 U3208 ( .A(n3160), .Q(n3143) );
  BUF15 U3209 ( .A(N2542), .Q(n3249) );
  INV4 U3210 ( .A(n3700), .Q(n3374) );
  BUF6 U3211 ( .A(n3565), .Q(n3290) );
  IMUX24 U3212 ( .A(net712307), .B(n3933), .S(n3932), .Q(n3934) );
  NAND28 U3213 ( .A(n3498), .B(n3499), .Q(net718339) );
  INV6 U3214 ( .A(n3828), .Q(n3499) );
  INV6 U3215 ( .A(n3027), .Q(n3037) );
  CLKIN6 U3216 ( .A(net712945), .Q(net715508) );
  INV4 U3217 ( .A(net712934), .Q(net712945) );
  NAND24 U3218 ( .A(net712167), .B(net725473), .Q(net712089) );
  CLKIN6 U3219 ( .A(n3674), .Q(n3426) );
  BUF15 U3220 ( .A(net723538), .Q(net723577) );
  NAND26 U3221 ( .A(net712698), .B(net715480), .Q(net712655) );
  INV6 U3222 ( .A(net712612), .Q(net712698) );
  NAND23 U3223 ( .A(net725419), .B(net712864), .Q(n3225) );
  NAND23 U3224 ( .A(net712484), .B(net724566), .Q(n3792) );
  NAND22 U3225 ( .A(net715746), .B(N2863), .Q(n4196) );
  INV10 U3226 ( .A(net719327), .Q(net718129) );
  INV10 U3227 ( .A(n4225), .Q(n3574) );
  CLKIN8 U3228 ( .A(n3377), .Q(n3378) );
  CLKIN12 U3229 ( .A(net713193), .Q(net713141) );
  NAND21 U3230 ( .A(net713052), .B(net713047), .Q(n3060) );
  INV8 U3231 ( .A(net712710), .Q(net712518) );
  INV4 U3232 ( .A(n3706), .Q(n2956) );
  NAND28 U3233 ( .A(n3640), .B(net715506), .Q(n3641) );
  CLKIN6 U3234 ( .A(n3645), .Q(n3636) );
  CLKIN15 U3235 ( .A(n3989), .Q(n4013) );
  NOR23 U3236 ( .A(n3475), .B(net712502), .Q(n3813) );
  NOR24 U3237 ( .A(n3474), .B(net718466), .Q(n3475) );
  NAND33 U3238 ( .A(net712089), .B(net726012), .C(n3283), .Q(n4225) );
  NAND26 U3239 ( .A(n2868), .B(n3101), .Q(n3099) );
  NAND23 U3240 ( .A(n2937), .B(n2938), .Q(net712672) );
  NAND23 U3241 ( .A(n3636), .B(n3635), .Q(net712893) );
  NAND32 U3242 ( .A(net723883), .B(net712722), .C(n3688), .Q(n3713) );
  XNR22 U3243 ( .A(net715608), .B(n3094), .Q(n3093) );
  NAND24 U3244 ( .A(net712803), .B(n3672), .Q(n3377) );
  CLKIN12 U3245 ( .A(net724932), .Q(n3169) );
  NAND22 U3246 ( .A(n3127), .B(net715616), .Q(net712729) );
  CLKIN6 U3247 ( .A(n2988), .Q(net713102) );
  INV4 U3248 ( .A(n2997), .Q(n2995) );
  NAND28 U3249 ( .A(net713142), .B(net713141), .Q(n3598) );
  OAI212 U3250 ( .A(arg[25]), .B(net713053), .C(n3613), .Q(n3615) );
  INV6 U3251 ( .A(net713053), .Q(net713104) );
  NAND22 U3252 ( .A(net724116), .B(net713053), .Q(n3072) );
  AOI312 U3253 ( .A(arg[25]), .B(net713055), .C(net713053), .D(n3612), .Q(
        n3613) );
  XNR22 U3254 ( .A(arg[26]), .B(net713096), .Q(n3601) );
  NAND24 U3255 ( .A(net724167), .B(net713196), .Q(net713100) );
  IMUX24 U3256 ( .A(N1905), .B(n3563), .S(n2959), .Q(net712113) );
  NAND24 U3257 ( .A(n3181), .B(n3163), .Q(n3160) );
  CLKIN6 U3258 ( .A(n3712), .Q(n3468) );
  CLKIN4 U3259 ( .A(net712934), .Q(net715510) );
  NAND26 U3260 ( .A(net712934), .B(net712976), .Q(net712980) );
  NOR33 U3261 ( .A(n3170), .B(n2961), .C(n3171), .Q(n3164) );
  INV12 U3262 ( .A(n3635), .Q(n3678) );
  OAI212 U3263 ( .A(net715450), .B(net712573), .C(net712655), .Q(n3162) );
  XNR22 U3264 ( .A(arg[26]), .B(net713096), .Q(net713143) );
  INV6 U3265 ( .A(net723547), .Q(net715678) );
  NAND28 U3266 ( .A(net712484), .B(n3818), .Q(n3789) );
  NOR22 U3267 ( .A(n2933), .B(N1786), .Q(n3957) );
  CLKIN8 U3268 ( .A(n4086), .Q(N2551) );
  IMUX22 U3269 ( .A(n3298), .B(N2488), .S(n2900), .Q(n4086) );
  NAND21 U3270 ( .A(n3679), .B(net725453), .Q(n3215) );
  NOR32 U3271 ( .A(n3279), .B(n3664), .C(n3665), .Q(n3648) );
  CLKIN6 U3272 ( .A(n3748), .Q(n3749) );
  INV6 U3273 ( .A(net723555), .Q(net712755) );
  NAND23 U3274 ( .A(n3091), .B(net712766), .Q(net712732) );
  OAI211 U3275 ( .A(net715768), .B(n3050), .C(net712903), .Q(n3045) );
  NAND26 U3276 ( .A(net712803), .B(n3652), .Q(net712864) );
  NAND22 U3277 ( .A(n3385), .B(n3386), .Q(n3759) );
  NAND26 U3278 ( .A(n3511), .B(n3512), .Q(n3858) );
  NAND26 U3279 ( .A(net712918), .B(net715678), .Q(n3645) );
  CLKIN12 U3280 ( .A(n3549), .Q(n3550) );
  NAND22 U3281 ( .A(n3998), .B(n4002), .Q(n3908) );
  NAND24 U3282 ( .A(net712145), .B(net715783), .Q(net718447) );
  INV6 U3283 ( .A(n3797), .Q(n3484) );
  NAND26 U3284 ( .A(n3812), .B(net725117), .Q(net712503) );
  NAND26 U3285 ( .A(net724188), .B(net724863), .Q(n3765) );
  NAND33 U3286 ( .A(net719152), .B(net715576), .C(n3653), .Q(n3488) );
  INV3 U3287 ( .A(n3930), .Q(n3833) );
  INV6 U3288 ( .A(N1782), .Q(n3974) );
  INV3 U3289 ( .A(net724863), .Q(n3183) );
  NOR21 U3290 ( .A(net721629), .B(net715776), .Q(n3391) );
  NAND26 U3291 ( .A(n3375), .B(n3376), .Q(n3762) );
  NAND26 U3292 ( .A(n3680), .B(net715705), .Q(n3681) );
  INV6 U3293 ( .A(n3681), .Q(n3455) );
  INV6 U3294 ( .A(net726138), .Q(net712020) );
  INV12 U3295 ( .A(n3543), .Q(n3935) );
  BUF2 U3296 ( .A(net723417), .Q(net726353) );
  NAND23 U3297 ( .A(n3208), .B(net725476), .Q(n3209) );
  INV2 U3298 ( .A(net717453), .Q(net721629) );
  NAND22 U3299 ( .A(net720041), .B(n3463), .Q(n3464) );
  NOR23 U3300 ( .A(net715610), .B(n3127), .Q(n3102) );
  INV6 U3301 ( .A(n4097), .Q(n4240) );
  INV8 U3302 ( .A(n4065), .Q(n4239) );
  INV3 U3303 ( .A(N2294), .Q(n4058) );
  NAND22 U3304 ( .A(net715480), .B(net712462), .Q(net712410) );
  NAND23 U3305 ( .A(net712589), .B(net715576), .Q(net712620) );
  XOR21 U3306 ( .A(net712970), .B(net715616), .Q(n3630) );
  NAND24 U3307 ( .A(net713120), .B(net713046), .Q(n2988) );
  INV1 U3308 ( .A(net715711), .Q(net725112) );
  CLKIN3 U3309 ( .A(net713130), .Q(net723480) );
  INV12 U3310 ( .A(net713090), .Q(net713087) );
  NAND23 U3311 ( .A(n4158), .B(n4157), .Q(n4285) );
  XNR21 U3312 ( .A(net723961), .B(n3859), .Q(n4000) );
  CLKBU12 U3313 ( .A(net712148), .Q(net715712) );
  NAND22 U3314 ( .A(n3230), .B(net712139), .Q(n4041) );
  INV8 U3315 ( .A(net710022), .Q(net713096) );
  NAND26 U3316 ( .A(n4033), .B(n4034), .Q(net718534) );
  INV6 U3317 ( .A(net717814), .Q(net715766) );
  CLKBU8 U3318 ( .A(net710022), .Q(net723547) );
  INV12 U3319 ( .A(arg[24]), .Q(net713055) );
  INV3 U3320 ( .A(net713146), .Q(n2996) );
  INV0 U3321 ( .A(n3866), .Q(n3399) );
  CLKIN12 U3322 ( .A(n4075), .Q(n4249) );
  INV12 U3323 ( .A(n4106), .Q(N2549) );
  XOR22 U3324 ( .A(net712782), .B(n3687), .Q(n2924) );
  INV8 U3325 ( .A(arg[25]), .Q(net713153) );
  INV3 U3326 ( .A(n3718), .Q(n3703) );
  INV10 U3327 ( .A(n3025), .Q(n3017) );
  NOR24 U3328 ( .A(arg[26]), .B(arg[27]), .Q(n3280) );
  INV8 U3329 ( .A(net703634), .Q(net715576) );
  CLKIN4 U3330 ( .A(net712935), .Q(net720967) );
  INV3 U3331 ( .A(net712879), .Q(n2947) );
  INV12 U3332 ( .A(net712938), .Q(n3034) );
  NAND28 U3333 ( .A(net724738), .B(net712963), .Q(n3063) );
  NAND28 U3334 ( .A(net718343), .B(net713072), .Q(net724738) );
  INV3 U3335 ( .A(net715510), .Q(net715506) );
  CLKIN15 U3336 ( .A(n3113), .Q(net712816) );
  CLKIN6 U3337 ( .A(n3688), .Q(n3222) );
  NAND26 U3338 ( .A(net712824), .B(net715680), .Q(n2944) );
  CLKIN12 U3339 ( .A(n3683), .Q(n3367) );
  INV4 U3340 ( .A(net712803), .Q(net712788) );
  CLKIN6 U3341 ( .A(n3835), .Q(n3234) );
  NAND28 U3342 ( .A(net712758), .B(net715572), .Q(net723768) );
  NAND22 U3343 ( .A(net723431), .B(net715678), .Q(n3881) );
  CLKIN1 U3344 ( .A(net715700), .Q(n2927) );
  OAI212 U3345 ( .A(net715450), .B(N1785), .C(net715711), .Q(n3978) );
  INV8 U3346 ( .A(net712133), .Q(net712132) );
  MUX26 U3347 ( .A(N2095), .B(n2894), .S(net712079), .Q(n2925) );
  MUX24 U3348 ( .A(N2109), .B(N1980), .S(n3578), .Q(n2926) );
  INV15 U3349 ( .A(net715719), .Q(net719234) );
  NAND28 U3350 ( .A(n3452), .B(n3453), .Q(n3454) );
  CLKIN3 U3351 ( .A(net715753), .Q(net720329) );
  INV6 U3352 ( .A(net719964), .Q(net722433) );
  CLKIN6 U3353 ( .A(net720329), .Q(net721034) );
  INV6 U3354 ( .A(n3136), .Q(N1777) );
  NAND24 U3355 ( .A(N2479), .B(net718128), .Q(n4094) );
  NAND26 U3356 ( .A(N2481), .B(net718128), .Q(n4091) );
  NAND24 U3357 ( .A(n3137), .B(net712434), .Q(net712433) );
  INV12 U3358 ( .A(net715646), .Q(net715642) );
  NAND26 U3359 ( .A(n3366), .B(n3367), .Q(net722205) );
  INV4 U3360 ( .A(n3702), .Q(n3686) );
  NAND21 U3361 ( .A(n3706), .B(net721083), .Q(n2957) );
  NAND28 U3362 ( .A(net712753), .B(net715608), .Q(n3688) );
  NAND26 U3363 ( .A(n3722), .B(net712825), .Q(net720699) );
  NAND23 U3364 ( .A(net715416), .B(arg[11]), .Q(n3194) );
  NAND21 U3365 ( .A(n3156), .B(net726353), .Q(n2930) );
  NAND24 U3366 ( .A(n2930), .B(n2931), .Q(n3142) );
  INV6 U3367 ( .A(net726353), .Q(n2929) );
  INV6 U3368 ( .A(n3142), .Q(n3176) );
  NAND23 U3369 ( .A(n4149), .B(n4150), .Q(n4270) );
  NAND23 U3370 ( .A(n4048), .B(net715768), .Q(net712147) );
  NOR32 U3371 ( .A(n3880), .B(n4004), .C(n3879), .Q(n2932) );
  INV3 U3372 ( .A(n2932), .Q(n2933) );
  INV1 U3373 ( .A(n4008), .Q(n3880) );
  INV6 U3374 ( .A(net723431), .Q(net712414) );
  NAND23 U3375 ( .A(N1922), .B(net725944), .Q(n4035) );
  NOR24 U3376 ( .A(N1917), .B(N1920), .Q(n4030) );
  CLKIN6 U3377 ( .A(net712644), .Q(n3101) );
  INV4 U3378 ( .A(net712942), .Q(n2963) );
  XNR20 U3379 ( .A(net721834), .B(n3738), .Q(n2935) );
  NAND24 U3380 ( .A(n3737), .B(net715540), .Q(n3738) );
  NAND24 U3381 ( .A(net724125), .B(n3634), .Q(n3404) );
  OAI211 U3382 ( .A(arg[26]), .B(net713157), .C(arg[27]), .Q(n3310) );
  OAI211 U3383 ( .A(net713097), .B(net713098), .C(n3310), .Q(n3603) );
  NAND22 U3384 ( .A(n3685), .B(net712790), .Q(n3447) );
  INV4 U3385 ( .A(n3685), .Q(n3446) );
  CLKIN0 U3386 ( .A(net715540), .Q(net722399) );
  CLKIN3 U3387 ( .A(net712910), .Q(net718388) );
  NAND22 U3388 ( .A(n3641), .B(net720185), .Q(n2938) );
  INV4 U3389 ( .A(n3641), .Q(n2936) );
  INV3 U3390 ( .A(net720185), .Q(n2951) );
  INV8 U3391 ( .A(net712967), .Q(net712865) );
  NAND33 U3392 ( .A(n2868), .B(net712688), .C(n2945), .Q(n3098) );
  INV2 U3393 ( .A(n3690), .Q(n2939) );
  INV3 U3394 ( .A(arg[27]), .Q(net713184) );
  NAND28 U3395 ( .A(n3468), .B(net718495), .Q(n3470) );
  NAND28 U3396 ( .A(net712731), .B(n3394), .Q(n3708) );
  NOR32 U3397 ( .A(n3708), .B(net712727), .C(net715680), .Q(n3711) );
  INV12 U3398 ( .A(n3708), .Q(n3714) );
  CLKIN3 U3399 ( .A(n3717), .Q(n3242) );
  NAND28 U3400 ( .A(n2940), .B(n2941), .Q(n2943) );
  NAND28 U3401 ( .A(n2942), .B(n2943), .Q(net712589) );
  CLKIN6 U3402 ( .A(n3134), .Q(n2940) );
  CLKIN3 U3403 ( .A(net712753), .Q(net723742) );
  INV3 U3404 ( .A(net723547), .Q(net715680) );
  INV3 U3405 ( .A(n3222), .Q(n2946) );
  NAND22 U3406 ( .A(net712879), .B(net712865), .Q(n2949) );
  NAND26 U3407 ( .A(n2947), .B(n2948), .Q(n2950) );
  NAND28 U3408 ( .A(n2949), .B(n2950), .Q(n3647) );
  CLKIN6 U3409 ( .A(net712865), .Q(n2948) );
  NOR24 U3410 ( .A(n3711), .B(n3710), .Q(n3459) );
  NAND28 U3411 ( .A(n3682), .B(n3378), .Q(n3673) );
  NAND24 U3412 ( .A(n3682), .B(net715704), .Q(n3683) );
  NAND20 U3413 ( .A(n2904), .B(net720697), .Q(n3775) );
  NAND26 U3414 ( .A(net712186), .B(net721410), .Q(net712184) );
  NAND28 U3415 ( .A(net712880), .B(n3467), .Q(n3246) );
  CLKIN15 U3416 ( .A(n3574), .Q(n3575) );
  NOR32 U3417 ( .A(net712721), .B(net715678), .C(n3222), .Q(n3223) );
  CLKIN12 U3418 ( .A(net712688), .Q(net712642) );
  NAND26 U3419 ( .A(net725420), .B(net723472), .Q(n3224) );
  NAND22 U3420 ( .A(net712164), .B(net712165), .Q(n3428) );
  NAND28 U3421 ( .A(net722204), .B(net722205), .Q(net721315) );
  NAND24 U3422 ( .A(n3681), .B(net723419), .Q(n3456) );
  INV6 U3423 ( .A(n3102), .Q(n3133) );
  IMUX24 U3424 ( .A(n3742), .B(n3741), .S(net721629), .Q(net712637) );
  NAND22 U3425 ( .A(n3464), .B(net715540), .Q(n3741) );
  CLKIN10 U3426 ( .A(net712733), .Q(net712821) );
  INV12 U3427 ( .A(n3656), .Q(n3401) );
  NAND22 U3428 ( .A(n3790), .B(net712536), .Q(n2953) );
  NAND24 U3429 ( .A(arg[15]), .B(n2952), .Q(n2954) );
  NAND24 U3430 ( .A(n2953), .B(n2954), .Q(n3843) );
  INV6 U3431 ( .A(net712536), .Q(n2952) );
  NAND23 U3432 ( .A(n3843), .B(net720783), .Q(n3940) );
  INV4 U3433 ( .A(n3843), .Q(n3208) );
  BUF2 U3434 ( .A(net712607), .Q(net720253) );
  INV6 U3435 ( .A(n3808), .Q(n3824) );
  CLKIN6 U3436 ( .A(net712864), .Q(net725420) );
  NAND28 U3437 ( .A(net712587), .B(net712588), .Q(net712462) );
  NAND26 U3438 ( .A(net712732), .B(n3692), .Q(n3693) );
  NAND23 U3439 ( .A(net712788), .B(arg[18]), .Q(n3449) );
  INV1 U3440 ( .A(net712781), .Q(net712727) );
  NAND28 U3441 ( .A(n3436), .B(net715576), .Q(net712781) );
  NAND24 U3442 ( .A(n2955), .B(n2956), .Q(n2958) );
  INV1 U3443 ( .A(net721083), .Q(n2955) );
  NAND22 U3444 ( .A(n3705), .B(net702066), .Q(n3706) );
  NAND23 U3445 ( .A(net712952), .B(net712935), .Q(net712951) );
  INV12 U3446 ( .A(N2063), .Q(n2959) );
  NAND28 U3447 ( .A(n3497), .B(n3618), .Q(n3296) );
  NOR24 U3448 ( .A(net720967), .B(net712966), .Q(n3409) );
  CLKIN6 U3449 ( .A(net712952), .Q(net712966) );
  NAND28 U3450 ( .A(n3362), .B(net722234), .Q(n3364) );
  NAND24 U3451 ( .A(net712946), .B(net718388), .Q(n3407) );
  INV15 U3452 ( .A(net703782), .Q(net715614) );
  XOR22 U3453 ( .A(net712980), .B(net712977), .Q(n2960) );
  INV12 U3454 ( .A(net712855), .Q(net712877) );
  NAND23 U3455 ( .A(net712885), .B(net715712), .Q(net712810) );
  NOR33 U3456 ( .A(net715572), .B(net712929), .C(net712816), .Q(n3120) );
  INV2 U3457 ( .A(net724932), .Q(n2961) );
  NAND22 U3458 ( .A(net712942), .B(n2876), .Q(n2964) );
  NAND24 U3459 ( .A(n2963), .B(n2962), .Q(n2965) );
  NAND26 U3460 ( .A(n2964), .B(n2965), .Q(net712804) );
  INV2 U3461 ( .A(n2876), .Q(n2962) );
  INV4 U3462 ( .A(net712804), .Q(net712888) );
  INV10 U3463 ( .A(n3626), .Q(n3411) );
  INV10 U3464 ( .A(n3080), .Q(net718604) );
  NAND22 U3465 ( .A(n3684), .B(n3683), .Q(net722204) );
  NAND28 U3466 ( .A(n3029), .B(net712991), .Q(n3056) );
  NAND28 U3467 ( .A(n3111), .B(n3112), .Q(net712803) );
  NAND22 U3468 ( .A(n3849), .B(n3821), .Q(n3852) );
  NAND24 U3469 ( .A(net712842), .B(net715608), .Q(n3123) );
  CLKIN6 U3470 ( .A(net712746), .Q(net712744) );
  NAND24 U3471 ( .A(net723742), .B(net715616), .Q(net712746) );
  NAND22 U3472 ( .A(net723637), .B(n3819), .Q(n3822) );
  NAND28 U3473 ( .A(n3077), .B(net720693), .Q(n3079) );
  NAND24 U3474 ( .A(net713112), .B(n3067), .Q(n3066) );
  NAND26 U3475 ( .A(n3088), .B(n3089), .Q(n3062) );
  NAND23 U3476 ( .A(net713141), .B(net713142), .Q(net713053) );
  AOI311 U3477 ( .A(net713143), .B(net713142), .C(net713141), .D(net715712), 
        .Q(n3071) );
  NAND21 U3478 ( .A(net713141), .B(net713142), .Q(net703634) );
  BUF12 U3479 ( .A(N2538), .Q(n3554) );
  CLKIN12 U3480 ( .A(net719237), .Q(net720894) );
  NAND22 U3481 ( .A(N2675), .B(net721268), .Q(n4110) );
  NAND26 U3482 ( .A(n2966), .B(net712323), .Q(n3138) );
  INV6 U3483 ( .A(n3248), .Q(n3891) );
  INV12 U3484 ( .A(n3657), .Q(n3674) );
  INV12 U3485 ( .A(n3137), .Q(net712211) );
  NAND24 U3486 ( .A(N2480), .B(net723620), .Q(n4092) );
  INV0 U3487 ( .A(net721315), .Q(net717806) );
  CLKIN6 U3488 ( .A(net712788), .Q(net718624) );
  NAND28 U3489 ( .A(n3785), .B(net715450), .Q(net712361) );
  NAND22 U3490 ( .A(net726021), .B(n3153), .Q(n3152) );
  NAND26 U3491 ( .A(n3796), .B(n3485), .Q(n3820) );
  NAND22 U3492 ( .A(n3518), .B(net722422), .Q(n3452) );
  MUX26 U3493 ( .A(n3523), .B(N2303), .S(net715717), .Q(n3518) );
  NAND26 U3494 ( .A(n3950), .B(net715614), .Q(n3836) );
  NAND22 U3495 ( .A(n3140), .B(n2901), .Q(n2966) );
  BUF12 U3496 ( .A(net712286), .Q(net715700) );
  INV0 U3497 ( .A(n2927), .Q(net724072) );
  NAND24 U3498 ( .A(n3945), .B(n3946), .Q(net712311) );
  INV15 U3499 ( .A(net712208), .Q(net715416) );
  NAND23 U3500 ( .A(net712145), .B(net715480), .Q(net712165) );
  INV6 U3501 ( .A(n4067), .Q(n4236) );
  CLKIN6 U3502 ( .A(net712732), .Q(net712716) );
  BUF15 U3503 ( .A(n4280), .Q(n3551) );
  NAND23 U3504 ( .A(N2484), .B(net723620), .Q(n2968) );
  NAND26 U3505 ( .A(net712934), .B(n3630), .Q(net712967) );
  NAND24 U3506 ( .A(net712521), .B(net712483), .Q(n3811) );
  IMUX24 U3507 ( .A(n4255), .B(N2306), .S(net715717), .Q(n4075) );
  INV6 U3508 ( .A(n4276), .Q(n3547) );
  INV3 U3509 ( .A(net716101), .Q(net726169) );
  NAND26 U3510 ( .A(net711940), .B(net711939), .Q(net703797) );
  CLKIN6 U3511 ( .A(n2972), .Q(n2973) );
  AOI312 U3512 ( .A(net725117), .B(n3976), .C(net723444), .D(n3975), .Q(n3981)
         );
  CLKIN6 U3513 ( .A(n3154), .Q(n3175) );
  OAI212 U3514 ( .A(net715788), .B(net712311), .C(net712286), .Q(net712307) );
  NOR42 U3515 ( .A(net712190), .B(net712189), .C(net712132), .D(net712131), 
        .Q(net712188) );
  CLKIN6 U3516 ( .A(net712165), .Q(net712189) );
  BUF6 U3517 ( .A(net713160), .Q(n2967) );
  CLKIN6 U3518 ( .A(n4034), .Q(N1977) );
  CLKIN3 U3519 ( .A(net712475), .Q(net723891) );
  NAND33 U3520 ( .A(net713150), .B(net713149), .C(net713151), .Q(n2994) );
  INV3 U3521 ( .A(net724429), .Q(net724923) );
  CLKIN3 U3522 ( .A(net724758), .Q(net725636) );
  CLKIN6 U3523 ( .A(n4061), .Q(n4244) );
  CLKIN3 U3524 ( .A(N2096), .Q(n3328) );
  INV3 U3525 ( .A(net716222), .Q(net723106) );
  CLKIN6 U3526 ( .A(n4052), .Q(n4252) );
  INV3 U3527 ( .A(n3022), .Q(n3023) );
  INV0 U3528 ( .A(n3350), .Q(n4116) );
  CLKIN6 U3529 ( .A(net716389), .Q(net716390) );
  INV12 U3530 ( .A(N1975), .Q(net712145) );
  INV3 U3531 ( .A(net712990), .Q(net719166) );
  NAND23 U3532 ( .A(n3085), .B(n3086), .Q(n3065) );
  NAND23 U3533 ( .A(N2870), .B(net719548), .Q(n4185) );
  XNR21 U3534 ( .A(n3797), .B(net712139), .Q(n3793) );
  NAND22 U3535 ( .A(n3484), .B(net724864), .Q(n3485) );
  NAND22 U3536 ( .A(net712976), .B(net712881), .Q(n3467) );
  CLKIN12 U3537 ( .A(n4093), .Q(n4291) );
  INV3 U3538 ( .A(net720783), .Q(net725476) );
  CLKIN3 U3539 ( .A(n3716), .Q(n3717) );
  INV3 U3540 ( .A(net715678), .Q(net725513) );
  NAND26 U3541 ( .A(net713011), .B(net713073), .Q(net712996) );
  INV3 U3542 ( .A(n3312), .Q(n3307) );
  CLKIN3 U3543 ( .A(n3237), .Q(n4068) );
  NAND24 U3544 ( .A(n3935), .B(n3388), .Q(n3946) );
  INV3 U3545 ( .A(n3419), .Q(n3420) );
  NAND26 U3546 ( .A(n3360), .B(n3361), .Q(n4010) );
  INV3 U3547 ( .A(net723881), .Q(net723927) );
  NAND22 U3548 ( .A(n3725), .B(net721162), .Q(n3732) );
  XNR21 U3549 ( .A(n3684), .B(n3367), .Q(n3725) );
  INV3 U3550 ( .A(net721162), .Q(net721834) );
  CLKIN12 U3551 ( .A(net712646), .Q(net712677) );
  INV1 U3552 ( .A(net712929), .Q(net723472) );
  INV3 U3553 ( .A(net713152), .Q(net713045) );
  INV3 U3554 ( .A(n4120), .Q(n3217) );
  INV12 U3555 ( .A(net712020), .Q(net660303) );
  CLKIN6 U3556 ( .A(net725635), .Q(n3139) );
  NAND26 U3557 ( .A(net723873), .B(net715788), .Q(net712501) );
  BUF2 U3558 ( .A(n3063), .Q(n3275) );
  INV3 U3559 ( .A(net724284), .Q(net712993) );
  INV3 U3560 ( .A(arg[23]), .Q(net713067) );
  XOR21 U3561 ( .A(n2897), .B(net713055), .Q(net724284) );
  NAND22 U3562 ( .A(net718618), .B(net718619), .Q(n3076) );
  NAND22 U3563 ( .A(net720826), .B(net713153), .Q(net718619) );
  XNR20 U3564 ( .A(arg[26]), .B(net713087), .Q(net713114) );
  INV3 U3565 ( .A(n3532), .Q(n3332) );
  INV3 U3566 ( .A(N2091), .Q(n3331) );
  INV3 U3567 ( .A(N1903), .Q(net721443) );
  NAND22 U3568 ( .A(n4005), .B(n4008), .Q(n3904) );
  NAND23 U3569 ( .A(net712702), .B(net715540), .Q(n3168) );
  INV3 U3570 ( .A(net712898), .Q(net722223) );
  INV3 U3571 ( .A(net721024), .Q(net722222) );
  CLKIN3 U3572 ( .A(net712899), .Q(n3049) );
  INV6 U3573 ( .A(n3076), .Q(net720693) );
  INV0 U3574 ( .A(net713127), .Q(net713078) );
  INV12 U3575 ( .A(arg[31]), .Q(net717816) );
  INV3 U3576 ( .A(n4206), .Q(n3405) );
  CLKIN1 U3577 ( .A(n3284), .Q(n3285) );
  IMUX23 U3578 ( .A(N1914), .B(n3396), .S(net715406), .Q(n4034) );
  NAND31 U3579 ( .A(net713170), .B(net713055), .C(net713153), .Q(n3005) );
  CLKIN3 U3580 ( .A(net715766), .Q(net715767) );
  NAND24 U3581 ( .A(n3320), .B(net723251), .Q(n3322) );
  NAND24 U3582 ( .A(net719964), .B(n3434), .Q(n3435) );
  INV3 U3583 ( .A(n4195), .Q(n3434) );
  NAND22 U3584 ( .A(n3433), .B(n3586), .Q(net712148) );
  NAND32 U3585 ( .A(net713189), .B(net719616), .C(net719953), .Q(n3433) );
  BUF6 U3586 ( .A(net712148), .Q(net715711) );
  BUF2 U3587 ( .A(net715540), .Q(net724566) );
  BUF2 U3588 ( .A(net724566), .Q(net720783) );
  INV3 U3589 ( .A(net715610), .Q(net715608) );
  BUF6 U3590 ( .A(net675324), .Q(net715480) );
  INV3 U3591 ( .A(N2963), .Q(n3286) );
  BUF15 U3592 ( .A(N2547), .Q(net716366) );
  OAI212 U3593 ( .A(net718129), .B(net712020), .C(n2968), .Q(N2547) );
  BUF15 U3594 ( .A(net715344), .Q(net723620) );
  BUF2 U3595 ( .A(net716366), .Q(net726276) );
  INV12 U3596 ( .A(N2819), .Q(net715378) );
  NAND22 U3597 ( .A(net715374), .B(N2857), .Q(net711886) );
  NAND21 U3598 ( .A(net715374), .B(N2856), .Q(net711884) );
  CLKIN4 U3599 ( .A(net715378), .Q(net720325) );
  OAI212 U3600 ( .A(net720325), .B(n2969), .C(net711886), .Q(res_4_) );
  IMUX20 U3601 ( .A(net715450), .B(n2971), .S(net722521), .Q(sqroot[15]) );
  INV15 U3602 ( .A(net717814), .Q(net715450) );
  INV2 U3603 ( .A(N2965), .Q(n2971) );
  CLKIN6 U3604 ( .A(n2970), .Q(net722521) );
  NAND28 U3605 ( .A(N2947), .B(roundup), .Q(n2970) );
  CLKIN15 U3606 ( .A(n2970), .Q(net711876) );
  NAND24 U3607 ( .A(N2674), .B(net718162), .Q(n2972) );
  BUF15 U3608 ( .A(N2627), .Q(net718162) );
  AOI212 U3609 ( .A(net721041), .B(net716332), .C(n2973), .Q(net716331) );
  INV8 U3610 ( .A(net716331), .Q(net640122) );
  CLKIN3 U3611 ( .A(net711990), .Q(net716332) );
  INV2 U3612 ( .A(N2545), .Q(net711990) );
  BUF2 U3613 ( .A(net640122), .Q(net721440) );
  IMUX22 U3614 ( .A(net725214), .B(N2289), .S(net718011), .Q(n2974) );
  MUX26 U3615 ( .A(N2097), .B(n2866), .S(net712079), .Q(net725214) );
  BUF15 U3616 ( .A(N2243), .Q(net718011) );
  BUF2 U3617 ( .A(net660309), .Q(net723292) );
  IMUX24 U3618 ( .A(n2977), .B(net724795), .S(net716206), .Q(net716268) );
  CLKIN6 U3619 ( .A(net703782), .Q(net715616) );
  OAI212 U3620 ( .A(n2978), .B(n2975), .C(n2976), .Q(net712192) );
  AOI211 U3621 ( .A(net715416), .B(net716390), .C(net715450), .Q(n2976) );
  NOR41 U3622 ( .A(net712132), .B(net712131), .C(net712169), .D(net712168), 
        .Q(net712167) );
  CLKIN6 U3623 ( .A(N1909), .Q(n2977) );
  XOR22 U3624 ( .A(net723959), .B(net712433), .Q(net724795) );
  NAND43 U3625 ( .A(n2979), .B(net726165), .C(net712166), .D(net712188), .Q(
        net712186) );
  AOI2112 U3626 ( .A(net712175), .B(net720783), .C(n2980), .D(net712202), .Q(
        n2979) );
  CLKIN4 U3627 ( .A(net722738), .Q(net712175) );
  NAND22 U3628 ( .A(net712113), .B(net715816), .Q(net712171) );
  IMUX22 U3629 ( .A(N1901), .B(arg[8]), .S(net715416), .Q(net712202) );
  AOI222 U3630 ( .A(net721443), .B(net715402), .C(net726168), .D(net726169), 
        .Q(net726165) );
  INV3 U3631 ( .A(net712197), .Q(net712166) );
  CLKIN6 U3632 ( .A(net712164), .Q(net712190) );
  NAND26 U3633 ( .A(net712114), .B(net725513), .Q(net712164) );
  NAND34 U3634 ( .A(net726012), .B(net712089), .C(n2981), .Q(net712087) );
  NOR24 U3635 ( .A(net712123), .B(n2885), .Q(n2981) );
  NAND28 U3636 ( .A(net712151), .B(net718535), .Q(net712123) );
  INV15 U3637 ( .A(net712087), .Q(net712079) );
  INV3 U3638 ( .A(n2982), .Q(n2985) );
  NAND22 U3639 ( .A(n2984), .B(n2983), .Q(n2982) );
  INV2 U3640 ( .A(net712146), .Q(n2984) );
  INV6 U3641 ( .A(net712147), .Q(net712146) );
  OAI221 U3642 ( .A(net715608), .B(net712196), .C(net715572), .D(net712203), 
        .Q(n2983) );
  INV15 U3643 ( .A(net713104), .Q(net715572) );
  IMUX24 U3644 ( .A(N1910), .B(N1781), .S(net715416), .Q(net712203) );
  INV1 U3645 ( .A(net712132), .Q(net721408) );
  INV2 U3646 ( .A(net712134), .Q(n2986) );
  NAND24 U3647 ( .A(net718447), .B(net712164), .Q(net712134) );
  IMUX22 U3648 ( .A(N2103), .B(N1974), .S(net712079), .Q(n2987) );
  CLKIN6 U3649 ( .A(net712114), .Q(N1974) );
  CLKIN0 U3650 ( .A(net660260), .Q(net724429) );
  OAI212 U3651 ( .A(net713103), .B(net713102), .C(net715769), .Q(n2991) );
  INV6 U3652 ( .A(n2989), .Q(net713103) );
  INV2 U3653 ( .A(net715766), .Q(net715769) );
  OAI212 U3654 ( .A(net713118), .B(net713117), .C(n2991), .Q(net713109) );
  CLKIN3 U3655 ( .A(net713102), .Q(net720951) );
  XOR31 U3656 ( .A(net725112), .B(net713127), .C(n3026), .Q(net713120) );
  NAND24 U3657 ( .A(net710022), .B(net724116), .Q(net713127) );
  XNR22 U3658 ( .A(n2992), .B(net713125), .Q(n3026) );
  NAND24 U3659 ( .A(n3018), .B(n3019), .Q(n2993) );
  NAND22 U3660 ( .A(n3025), .B(arg[26]), .Q(n3018) );
  NAND28 U3661 ( .A(net722414), .B(net716402), .Q(n3025) );
  NAND26 U3662 ( .A(n3017), .B(net718490), .Q(n3019) );
  INV3 U3663 ( .A(arg[26]), .Q(net718490) );
  NAND24 U3664 ( .A(net713084), .B(net713085), .Q(net713125) );
  INV6 U3665 ( .A(net713121), .Q(net713046) );
  AOI212 U3666 ( .A(n2988), .B(n2989), .C(net715766), .Q(net725046) );
  NOR33 U3667 ( .A(n3021), .B(n2994), .C(n2995), .Q(net713121) );
  NAND23 U3668 ( .A(net713046), .B(net713045), .Q(net713044) );
  NAND24 U3669 ( .A(net713146), .B(net713148), .Q(n3021) );
  NAND28 U3670 ( .A(net713159), .B(n2967), .Q(net713148) );
  NAND22 U3671 ( .A(net713121), .B(arg[24]), .Q(net713052) );
  NAND23 U3672 ( .A(net713121), .B(net713130), .Q(n2989) );
  OAI222 U3673 ( .A(n3002), .B(n3001), .C(n3017), .D(net718490), .Q(n2997) );
  NOR42 U3674 ( .A(n2996), .B(net713138), .C(n2994), .D(n2995), .Q(net713031)
         );
  AOI2112 U3675 ( .A(n2990), .B(net715767), .C(n3003), .D(net713157), .Q(n3002) );
  OAI212 U3676 ( .A(n3024), .B(n3004), .C(n3005), .Q(n3003) );
  NOR21 U3677 ( .A(arg[26]), .B(arg[27]), .Q(n3024) );
  INV8 U3678 ( .A(net713129), .Q(net713157) );
  AOI2111 U3679 ( .A(net723527), .B(net713184), .C(n3007), .D(n3025), .Q(n3001) );
  OAI211 U3680 ( .A(net715450), .B(net713186), .C(n3005), .Q(n3007) );
  OAI212 U3681 ( .A(arg[28]), .B(net713197), .C(net723781), .Q(net713186) );
  NAND34 U3682 ( .A(n2997), .B(net713146), .C(net713148), .Q(net713158) );
  OAI212 U3683 ( .A(n3008), .B(n3009), .C(n3000), .Q(n3006) );
  NAND22 U3684 ( .A(n2990), .B(net710022), .Q(net713099) );
  CLKIN3 U3685 ( .A(net713211), .Q(n3008) );
  NOR23 U3686 ( .A(net720403), .B(n3011), .Q(n3009) );
  NAND26 U3687 ( .A(n2998), .B(n3023), .Q(n3000) );
  NAND31 U3688 ( .A(n3006), .B(net715450), .C(net713100), .Q(net713150) );
  CLKIN6 U3689 ( .A(n3011), .Q(n2998) );
  NAND21 U3690 ( .A(n3010), .B(net713199), .Q(n3022) );
  OAI212 U3691 ( .A(arg[27]), .B(arg[26]), .C(net719615), .Q(n3010) );
  INV15 U3692 ( .A(arg[28]), .Q(net719615) );
  NAND28 U3693 ( .A(n3020), .B(arg[30]), .Q(net713199) );
  INV2 U3694 ( .A(n3000), .Q(net713162) );
  OAI212 U3695 ( .A(n3008), .B(n3009), .C(n3000), .Q(net724021) );
  INV6 U3696 ( .A(n3012), .Q(n3011) );
  NAND22 U3697 ( .A(n2998), .B(net713167), .Q(net713166) );
  OAI2112 U3698 ( .A(n3014), .B(n3013), .C(n3015), .D(n3016), .Q(n3012) );
  NOR24 U3699 ( .A(arg[29]), .B(arg[30]), .Q(n3014) );
  OAI212 U3700 ( .A(arg[31]), .B(n2999), .C(net713171), .Q(n3013) );
  INV12 U3701 ( .A(arg[30]), .Q(n2999) );
  INV15 U3702 ( .A(arg[28]), .Q(net713171) );
  NAND33 U3703 ( .A(n3020), .B(arg[28]), .C(arg[30]), .Q(n3015) );
  INV15 U3704 ( .A(arg[31]), .Q(n3020) );
  NOR24 U3705 ( .A(arg[27]), .B(arg[26]), .Q(n3016) );
  AOI212 U3706 ( .A(n3030), .B(n3031), .C(n3037), .Q(net712942) );
  AOI211 U3707 ( .A(n3028), .B(net715710), .C(n3035), .Q(n3030) );
  INV6 U3708 ( .A(net712946), .Q(n3028) );
  BUF2 U3709 ( .A(net712148), .Q(net715710) );
  OAI222 U3710 ( .A(n3028), .B(n3036), .C(net715710), .D(net712950), .Q(n3035)
         );
  NAND22 U3711 ( .A(n3034), .B(net715480), .Q(n3036) );
  INV6 U3712 ( .A(net712950), .Q(net712914) );
  AOI312 U3713 ( .A(net715480), .B(net712946), .C(n3032), .D(n3033), .Q(n3031)
         );
  NAND28 U3714 ( .A(net712957), .B(net715825), .Q(net712946) );
  INV6 U3715 ( .A(net712951), .Q(n3032) );
  NOR42 U3716 ( .A(net715480), .B(n3032), .C(net712914), .D(n3034), .Q(n3033)
         );
  NAND24 U3717 ( .A(n3038), .B(n3039), .Q(n3027) );
  NOR23 U3718 ( .A(net712965), .B(n3037), .Q(net712960) );
  AOI2112 U3719 ( .A(n3042), .B(n3043), .C(net712894), .D(n3044), .Q(n3038) );
  AOI222 U3720 ( .A(net712983), .B(net712984), .C(net712985), .D(net716699), 
        .Q(n3039) );
  NOR24 U3721 ( .A(net715825), .B(net712957), .Q(net712983) );
  NOR24 U3722 ( .A(net712895), .B(net712910), .Q(net712984) );
  CLKIN3 U3723 ( .A(net719165), .Q(net712985) );
  OAI212 U3724 ( .A(net715572), .B(net712966), .C(n3027), .Q(net712959) );
  AOI212 U3725 ( .A(n3054), .B(n3055), .C(n3056), .Q(n3042) );
  NAND23 U3726 ( .A(n3062), .B(net715576), .Q(n3054) );
  NAND24 U3727 ( .A(net713067), .B(n3087), .Q(n3088) );
  NAND24 U3728 ( .A(arg[23]), .B(n3063), .Q(n3089) );
  NAND24 U3729 ( .A(n3061), .B(net712935), .Q(n3055) );
  NAND24 U3730 ( .A(net712940), .B(net712939), .Q(n3061) );
  NAND22 U3731 ( .A(net712970), .B(net712963), .Q(net712940) );
  NAND28 U3732 ( .A(arg[22]), .B(net715614), .Q(net712939) );
  NAND28 U3733 ( .A(n3057), .B(net715480), .Q(n3029) );
  NAND28 U3734 ( .A(net712992), .B(net715768), .Q(net712991) );
  NAND24 U3735 ( .A(n3051), .B(net715824), .Q(n3043) );
  XNR22 U3736 ( .A(n3052), .B(net724284), .Q(n3051) );
  XOR22 U3737 ( .A(net715576), .B(n3053), .Q(net712997) );
  BUF2 U3738 ( .A(net715674), .Q(net715824) );
  XNR22 U3739 ( .A(net713001), .B(net713002), .Q(net712894) );
  OAI2112 U3740 ( .A(n3045), .B(n3046), .C(net712898), .D(n3047), .Q(n3044) );
  CLKIN3 U3741 ( .A(net713024), .Q(n3050) );
  NAND23 U3742 ( .A(net720951), .B(net721341), .Q(net712903) );
  NAND22 U3743 ( .A(net713008), .B(n3050), .Q(net712902) );
  NAND26 U3744 ( .A(net713015), .B(net715450), .Q(net712898) );
  NAND22 U3745 ( .A(n3048), .B(n3049), .Q(n3047) );
  CLKIN0 U3746 ( .A(net712903), .Q(n3048) );
  NAND31 U3747 ( .A(net713020), .B(net713009), .C(net715767), .Q(net712899) );
  NAND26 U3748 ( .A(n3038), .B(net723514), .Q(net712934) );
  NAND28 U3749 ( .A(n3078), .B(n3079), .Q(n3057) );
  NAND22 U3750 ( .A(n3040), .B(n3076), .Q(n3078) );
  INV6 U3751 ( .A(n3058), .Q(n3040) );
  CLKIN6 U3752 ( .A(n3040), .Q(n3077) );
  OAI212 U3753 ( .A(net712904), .B(n3080), .C(n3059), .Q(n3058) );
  NAND26 U3754 ( .A(net713011), .B(net713073), .Q(net712904) );
  BUF15 U3755 ( .A(n3041), .Q(n3080) );
  XNR21 U3756 ( .A(net715674), .B(n3060), .Q(n3059) );
  INV1 U3757 ( .A(net715678), .Q(net715674) );
  NAND21 U3758 ( .A(n3053), .B(net713055), .Q(net713047) );
  CLKIN2 U3759 ( .A(n3040), .Q(net721548) );
  OAI222 U3760 ( .A(net713109), .B(n3064), .C(n3066), .D(n3065), .Q(n3041) );
  AOI312 U3761 ( .A(net713058), .B(net715711), .C(net724065), .D(n3074), .Q(
        n3064) );
  NAND24 U3762 ( .A(n3083), .B(n3084), .Q(n3074) );
  NAND26 U3763 ( .A(net713116), .B(net713045), .Q(n3075) );
  INV3 U3764 ( .A(net713043), .Q(n3081) );
  NAND22 U3765 ( .A(net723547), .B(net713153), .Q(net713043) );
  AOI222 U3766 ( .A(n3072), .B(n3071), .C(n3073), .D(net713052), .Q(net713117)
         );
  XOR22 U3767 ( .A(arg[26]), .B(net713087), .Q(net724116) );
  OAI210 U3768 ( .A(arg[22]), .B(n3053), .C(net713055), .Q(n3073) );
  NAND22 U3769 ( .A(net713067), .B(net712963), .Q(n3053) );
  NOR33 U3770 ( .A(net715480), .B(n3069), .C(n3070), .Q(net713118) );
  CLKIN12 U3771 ( .A(net713057), .Q(n3069) );
  CLKIN6 U3772 ( .A(net725046), .Q(net713112) );
  OAI221 U3773 ( .A(net723547), .B(net713114), .C(net723547), .D(net715480), 
        .Q(n3067) );
  NAND22 U3774 ( .A(arg[25]), .B(net713061), .Q(n3085) );
  INV6 U3775 ( .A(n3068), .Q(net713061) );
  NAND23 U3776 ( .A(net713153), .B(n3068), .Q(n3086) );
  NAND26 U3777 ( .A(net713116), .B(net713055), .Q(n3068) );
  OAI212 U3778 ( .A(net712904), .B(n3080), .C(net712963), .Q(net713068) );
  CLKIN0 U3779 ( .A(net712758), .Q(net723417) );
  BUF2 U3780 ( .A(net723742), .Q(n3134) );
  NAND26 U3781 ( .A(net702066), .B(n3093), .Q(n3092) );
  NAND26 U3782 ( .A(n3091), .B(n3135), .Q(net702066) );
  NAND22 U3783 ( .A(net712731), .B(net712730), .Q(n3094) );
  NAND24 U3784 ( .A(net721808), .B(net712743), .Q(net712731) );
  AOI212 U3785 ( .A(n3095), .B(net724789), .C(n3096), .Q(n3091) );
  OAI212 U3786 ( .A(net723702), .B(net712773), .C(net712774), .Q(n3135) );
  OAI2112 U3787 ( .A(net712784), .B(net712754), .C(net712746), .D(net712781), 
        .Q(net712773) );
  NOR42 U3788 ( .A(net724008), .B(net712777), .C(net712775), .D(net712778), 
        .Q(net712774) );
  NOR24 U3789 ( .A(n3130), .B(n3103), .Q(n3095) );
  CLKIN6 U3790 ( .A(n3129), .Q(n3130) );
  NOR24 U3791 ( .A(net724008), .B(n3132), .Q(n3129) );
  NAND28 U3792 ( .A(n3133), .B(net723883), .Q(n3132) );
  INV2 U3793 ( .A(net703782), .Q(net715610) );
  XNR22 U3794 ( .A(n3131), .B(n3108), .Q(n3127) );
  NAND28 U3795 ( .A(net724837), .B(net725513), .Q(net723883) );
  NAND33 U3796 ( .A(n3105), .B(n3104), .C(net712787), .Q(n3103) );
  NOR24 U3797 ( .A(net712642), .B(net712760), .Q(n3105) );
  INV3 U3798 ( .A(arg[16]), .Q(net712760) );
  XNR22 U3799 ( .A(n3106), .B(n3107), .Q(n3104) );
  OAI210 U3800 ( .A(net723435), .B(net712790), .C(net715788), .Q(n3106) );
  INV12 U3801 ( .A(net715508), .Q(net723435) );
  INV3 U3802 ( .A(arg[19]), .Q(net712790) );
  NAND22 U3803 ( .A(net723603), .B(net715788), .Q(n3107) );
  NAND22 U3804 ( .A(arg[18]), .B(net715705), .Q(net712787) );
  NAND43 U3805 ( .A(n3099), .B(n3098), .C(n3097), .D(n3100), .Q(n3096) );
  NAND28 U3806 ( .A(net712821), .B(net715711), .Q(net712644) );
  XNR22 U3807 ( .A(net723472), .B(net712864), .Q(net712824) );
  NAND26 U3808 ( .A(net712733), .B(net715480), .Q(net712688) );
  AOI2112 U3809 ( .A(net717453), .B(net715450), .C(net721379), .D(n3090), .Q(
        n3097) );
  CLKIN6 U3810 ( .A(net721166), .Q(net717453) );
  CLKIN12 U3811 ( .A(net712668), .Q(n3090) );
  NAND28 U3812 ( .A(net720699), .B(net720700), .Q(net712668) );
  NOR24 U3813 ( .A(net712677), .B(net721315), .Q(n3100) );
  BUF2 U3814 ( .A(net712860), .Q(n3131) );
  NAND28 U3815 ( .A(n3111), .B(n3112), .Q(net712792) );
  XNR21 U3816 ( .A(n3110), .B(net723435), .Q(n3109) );
  INV3 U3817 ( .A(net712881), .Q(n3110) );
  NAND22 U3818 ( .A(net712790), .B(net712793), .Q(net712881) );
  XNR22 U3819 ( .A(n3131), .B(n3108), .Q(net712752) );
  INV6 U3820 ( .A(n3115), .Q(n3111) );
  NOR24 U3821 ( .A(net712887), .B(n3114), .Q(n3112) );
  OAI312 U3822 ( .A(n3117), .B(n3118), .C(n3116), .D(n3119), .Q(n3115) );
  OAI211 U3823 ( .A(net715576), .B(n3121), .C(n3113), .Q(n3117) );
  XNR22 U3824 ( .A(net712879), .B(net712967), .Q(n3121) );
  NAND28 U3825 ( .A(net712848), .B(net725513), .Q(n3113) );
  AOI2112 U3826 ( .A(n3122), .B(n3123), .C(net712877), .D(n3124), .Q(n3116) );
  NAND28 U3827 ( .A(net712860), .B(net723435), .Q(net712880) );
  XNR22 U3828 ( .A(arg[21]), .B(net712979), .Q(net712842) );
  AOI212 U3829 ( .A(n3125), .B(net715608), .C(n3126), .Q(n3124) );
  AOI221 U3830 ( .A(net712945), .B(arg[21]), .C(net715508), .D(net712977), .Q(
        n3125) );
  CLKIN3 U3831 ( .A(arg[21]), .Q(net712977) );
  OAI212 U3832 ( .A(arg[18]), .B(net712881), .C(net712976), .Q(n3126) );
  CLKIN3 U3833 ( .A(arg[20]), .Q(net712976) );
  NAND22 U3834 ( .A(net712919), .B(net712815), .Q(n3118) );
  NAND26 U3835 ( .A(net715480), .B(net712917), .Q(net712815) );
  AOI312 U3836 ( .A(net712815), .B(net712919), .C(n3120), .D(n3128), .Q(n3119)
         );
  CLKIN6 U3837 ( .A(n3121), .Q(net712929) );
  NOR24 U3838 ( .A(net712810), .B(net712831), .Q(n3128) );
  NOR20 U3839 ( .A(net712831), .B(net712810), .Q(net721242) );
  OAI2112 U3840 ( .A(net712831), .B(net712893), .C(net712672), .D(net712674), 
        .Q(n3114) );
  XNR22 U3841 ( .A(net712330), .B(n3138), .Q(n3136) );
  INV3 U3842 ( .A(arg[13]), .Q(net712330) );
  NAND28 U3843 ( .A(n3140), .B(n2901), .Q(n3137) );
  CLKIN3 U3844 ( .A(arg[12]), .Q(net712323) );
  XNR22 U3845 ( .A(net712330), .B(n3138), .Q(net721714) );
  INV6 U3846 ( .A(n3144), .Q(n3140) );
  OAI212 U3847 ( .A(net712341), .B(n3145), .C(n3146), .Q(n3144) );
  INV6 U3848 ( .A(net712359), .Q(net712341) );
  NOR24 U3849 ( .A(n3155), .B(n3177), .Q(n3145) );
  INV2 U3850 ( .A(net712412), .Q(n3155) );
  NAND24 U3851 ( .A(net712369), .B(net715711), .Q(net712412) );
  NOR33 U3852 ( .A(n3175), .B(net715824), .C(n3176), .Q(n3177) );
  NAND23 U3853 ( .A(net712462), .B(net715480), .Q(n3154) );
  NOR42 U3854 ( .A(n3148), .B(net712216), .C(n2892), .D(n3147), .Q(n3146) );
  INV1 U3855 ( .A(net712415), .Q(n3148) );
  XNR22 U3856 ( .A(net712652), .B(net712656), .Q(net712415) );
  AOI212 U3857 ( .A(net712363), .B(n3139), .C(n3150), .Q(n3149) );
  NOR24 U3858 ( .A(net725636), .B(net723637), .Q(net725635) );
  OAI222 U3859 ( .A(n3151), .B(n3152), .C(net712357), .D(net712366), .Q(n3150)
         );
  INV6 U3860 ( .A(net712366), .Q(n3151) );
  CLKIN3 U3861 ( .A(net712560), .Q(n3153) );
  NAND28 U3862 ( .A(net712637), .B(net720124), .Q(net712357) );
  INV6 U3863 ( .A(net712544), .Q(net712238) );
  NAND28 U3864 ( .A(n3140), .B(n3141), .Q(net712286) );
  OAI212 U3865 ( .A(n3142), .B(net715680), .C(net712410), .Q(net712461) );
  XNR22 U3866 ( .A(net715576), .B(n3158), .Q(n3157) );
  NOR22 U3867 ( .A(net712596), .B(n3179), .Q(n3158) );
  NOR32 U3868 ( .A(n3183), .B(net712582), .C(n3178), .Q(n3179) );
  NAND28 U3869 ( .A(net724864), .B(net712503), .Q(net724863) );
  INV3 U3870 ( .A(net724188), .Q(n3178) );
  NAND43 U3871 ( .A(net712505), .B(net712504), .C(net712512), .D(net712503), 
        .Q(net724188) );
  INV15 U3872 ( .A(net706857), .Q(net715646) );
  CLKBU15 U3873 ( .A(net715642), .Q(net715816) );
  NAND28 U3874 ( .A(n3143), .B(net712529), .Q(net706857) );
  NOR23 U3875 ( .A(net723918), .B(net715646), .Q(net723917) );
  XNR22 U3876 ( .A(arg[14]), .B(net715646), .Q(net712316) );
  INV12 U3877 ( .A(net712600), .Q(net712529) );
  NAND26 U3878 ( .A(net706857), .B(net712454), .Q(net712536) );
  NAND23 U3879 ( .A(net712484), .B(net712478), .Q(net712496) );
  NAND26 U3880 ( .A(n3180), .B(n3182), .Q(n3181) );
  INV6 U3881 ( .A(n3161), .Q(n3180) );
  OAI2112 U3882 ( .A(net712610), .B(net712501), .C(n3173), .D(n3174), .Q(n3161) );
  INV2 U3883 ( .A(net712620), .Q(net712610) );
  OAI211 U3884 ( .A(net712507), .B(net712504), .C(net712620), .Q(n3173) );
  INV6 U3885 ( .A(net712513), .Q(net712507) );
  OAI212 U3886 ( .A(net715544), .B(net712760), .C(net712531), .Q(net712504) );
  OAI212 U3887 ( .A(n3169), .B(net712607), .C(net712620), .Q(n3174) );
  NOR23 U3888 ( .A(net712619), .B(n3162), .Q(n3182) );
  OAI312 U3889 ( .A(net712596), .B(n3164), .C(n3165), .D(n3166), .Q(n3163) );
  AOI312 U3890 ( .A(n3172), .B(net715544), .C(net723890), .D(n3159), .Q(n3171)
         );
  OAI210 U3891 ( .A(net712139), .B(net712712), .C(n2872), .Q(n3172) );
  INV3 U3892 ( .A(arg[17]), .Q(net712712) );
  INV6 U3893 ( .A(net702066), .Q(net715544) );
  XNR22 U3894 ( .A(arg[16]), .B(net715542), .Q(net723890) );
  INV6 U3895 ( .A(net712512), .Q(n3159) );
  NAND28 U3896 ( .A(net712518), .B(net712139), .Q(net712512) );
  AOI2112 U3897 ( .A(n3167), .B(net715608), .C(net715788), .D(n3184), .Q(n3165) );
  XOR22 U3898 ( .A(net718432), .B(n3168), .Q(n3167) );
  INV2 U3899 ( .A(net712700), .Q(net718432) );
  XNR21 U3900 ( .A(net725117), .B(net712755), .Q(net712702) );
  INV15 U3901 ( .A(net715542), .Q(net715540) );
  CLKIN6 U3902 ( .A(net723541), .Q(n3184) );
  INV2 U3903 ( .A(net723873), .Q(net723541) );
  NOR42 U3904 ( .A(net712607), .B(net723538), .C(net712555), .D(net712619), 
        .Q(n3166) );
  NOR24 U3905 ( .A(net719727), .B(net712612), .Q(net723538) );
  NAND24 U3906 ( .A(n3143), .B(net712529), .Q(net712521) );
  NAND28 U3907 ( .A(n3143), .B(net712529), .Q(net712484) );
  NAND28 U3908 ( .A(n3820), .B(net715788), .Q(n3821) );
  NAND20 U3909 ( .A(n3485), .B(net723435), .Q(n3185) );
  INV3 U3910 ( .A(n3185), .Q(n3186) );
  NAND22 U3911 ( .A(N2493), .B(net719306), .Q(n4080) );
  BUF2 U3912 ( .A(n3551), .Q(n3187) );
  CLKIN0 U3913 ( .A(n3548), .Q(n4193) );
  BUF12 U3914 ( .A(N2552), .Q(n3540) );
  AOI211 U3915 ( .A(net721041), .B(net726276), .C(n3557), .Q(n3278) );
  NAND24 U3916 ( .A(n4135), .B(n4136), .Q(n4263) );
  CLKIN6 U3917 ( .A(n4073), .Q(n4063) );
  IMUX22 U3918 ( .A(n4252), .B(N2298), .S(net715719), .Q(n4084) );
  CLKIN4 U3919 ( .A(N2288), .Q(n4062) );
  INV6 U3920 ( .A(N1971), .Q(n3341) );
  NAND24 U3921 ( .A(n4144), .B(n4143), .Q(n4217) );
  NAND23 U3922 ( .A(n4143), .B(n4144), .Q(n4267) );
  NAND21 U3923 ( .A(N2554), .B(net719447), .Q(n4144) );
  NAND22 U3924 ( .A(N2672), .B(net718162), .Q(n4113) );
  CLKIN6 U3925 ( .A(n3574), .Q(n3576) );
  NAND24 U3926 ( .A(n3264), .B(net719234), .Q(n3188) );
  NAND22 U3927 ( .A(N2292), .B(net715719), .Q(n3189) );
  NAND26 U3928 ( .A(n3188), .B(n3189), .Q(net726138) );
  INV8 U3929 ( .A(n3330), .Q(n4293) );
  CLKIN3 U3930 ( .A(net712199), .Q(net726092) );
  NAND24 U3931 ( .A(N1912), .B(net726092), .Q(n3190) );
  NAND28 U3932 ( .A(n3190), .B(n3191), .Q(N1975) );
  CLKIN12 U3933 ( .A(net722560), .Q(net722561) );
  BUF15 U3934 ( .A(n3273), .Q(n3192) );
  INV6 U3935 ( .A(net715739), .Q(net715360) );
  BUF2 U3936 ( .A(n4012), .Q(n3338) );
  BUF2 U3937 ( .A(net715416), .Q(net715412) );
  NAND23 U3938 ( .A(N2485), .B(net718129), .Q(n4088) );
  NAND28 U3939 ( .A(n3193), .B(n3194), .Q(net722729) );
  NAND24 U3940 ( .A(net712203), .B(net715572), .Q(net712133) );
  NOR22 U3941 ( .A(n3529), .B(net715544), .Q(n3565) );
  INV8 U3942 ( .A(n4099), .Q(n4238) );
  INV6 U3943 ( .A(n4015), .Q(N1979) );
  NAND24 U3944 ( .A(n3930), .B(n3929), .Q(n3845) );
  INV3 U3945 ( .A(n3995), .Q(n3992) );
  NAND41 U3946 ( .A(n2889), .B(n3997), .C(n3998), .D(n3991), .Q(n3995) );
  INV6 U3947 ( .A(n4066), .Q(n4237) );
  NAND24 U3948 ( .A(N1904), .B(net725903), .Q(n3193) );
  OAI310 U3949 ( .A(n3777), .B(net715544), .C(n3776), .D(n3775), .Q(n3782) );
  NAND20 U3950 ( .A(n3886), .B(net715678), .Q(n3838) );
  INV6 U3951 ( .A(n3886), .Q(n3864) );
  IMUX23 U3952 ( .A(N1908), .B(N1779), .S(net712199), .Q(n4039) );
  INV6 U3953 ( .A(n4049), .Q(n4255) );
  NAND26 U3954 ( .A(n3566), .B(net712139), .Q(n3929) );
  INV2 U3955 ( .A(n3929), .Q(n3847) );
  NAND21 U3956 ( .A(n3791), .B(n3792), .Q(n3197) );
  NAND24 U3957 ( .A(n3195), .B(n3196), .Q(n3198) );
  CLKIN3 U3958 ( .A(n3791), .Q(n3195) );
  CLKIN15 U3959 ( .A(net715348), .Q(net715344) );
  CLKIN8 U3960 ( .A(net715348), .Q(net715346) );
  CLKIN3 U3961 ( .A(n3977), .Q(n3199) );
  CLKIN6 U3962 ( .A(n3977), .Q(n3968) );
  INV2 U3963 ( .A(net712888), .Q(net723419) );
  NAND28 U3964 ( .A(net712789), .B(net725117), .Q(net712730) );
  INV1 U3965 ( .A(net712674), .Q(net712825) );
  BUF2 U3966 ( .A(n3341), .Q(n3200) );
  NAND24 U3967 ( .A(n3303), .B(net722422), .Q(n3201) );
  NAND22 U3968 ( .A(N2476), .B(net717907), .Q(n3202) );
  NAND28 U3969 ( .A(n3201), .B(n3202), .Q(n3400) );
  BUF15 U3970 ( .A(N2243), .Q(net715719) );
  NAND23 U3971 ( .A(n4156), .B(n4155), .Q(n4279) );
  INV4 U3972 ( .A(n4082), .Q(N2554) );
  INV8 U3973 ( .A(n4084), .Q(n4245) );
  BUF15 U3974 ( .A(N2541), .Q(n3203) );
  INV2 U3975 ( .A(net718067), .Q(net715725) );
  CLKIN12 U3976 ( .A(net715326), .Q(net719237) );
  INV4 U3977 ( .A(N2295), .Q(n4056) );
  INV8 U3978 ( .A(n3235), .Q(N2544) );
  NAND26 U3979 ( .A(n3323), .B(net722422), .Q(n3348) );
  NAND24 U3980 ( .A(n3856), .B(net715572), .Q(n3837) );
  BUF2 U3981 ( .A(net715704), .Q(net725733) );
  XOR21 U3982 ( .A(net712363), .B(n3902), .Q(n3515) );
  BUF2 U3983 ( .A(net712668), .Q(net721373) );
  CLKBU4 U3984 ( .A(n3760), .Q(n3410) );
  NAND21 U3985 ( .A(n3760), .B(net715678), .Q(n3385) );
  INV3 U3986 ( .A(n4038), .Q(n4040) );
  NAND24 U3987 ( .A(n4039), .B(net715788), .Q(n4038) );
  NAND26 U3988 ( .A(n3329), .B(n4088), .Q(N2548) );
  NAND26 U3989 ( .A(n3478), .B(net723912), .Q(n3479) );
  INV6 U3990 ( .A(n3777), .Q(n3734) );
  NAND22 U3991 ( .A(n3700), .B(n3288), .Q(n3375) );
  NAND24 U3992 ( .A(n3662), .B(net712792), .Q(n3663) );
  INV3 U3993 ( .A(n3739), .Q(n3740) );
  CLKIN1 U3994 ( .A(net712529), .Q(net721638) );
  CLKIN6 U3995 ( .A(net722422), .Q(net725641) );
  INV0 U3996 ( .A(n3820), .Q(n3932) );
  INV15 U3997 ( .A(net718324), .Q(net719306) );
  CLKBU15 U3998 ( .A(net719293), .Q(net718226) );
  NAND20 U3999 ( .A(n3229), .B(net718324), .Q(n3503) );
  NAND23 U4000 ( .A(net720325), .B(N2859), .Q(n4202) );
  CLKIN4 U4001 ( .A(net720325), .Q(net719964) );
  NAND22 U4002 ( .A(N2678), .B(net721268), .Q(n4105) );
  CLKIN6 U4003 ( .A(net721268), .Q(net722560) );
  NAND24 U4004 ( .A(n4142), .B(n4141), .Q(n4266) );
  BUF12 U4005 ( .A(N2627), .Q(net721268) );
  AOI211 U4006 ( .A(n3234), .B(n3849), .C(n3848), .Q(n3850) );
  MUX22 U4007 ( .A(n3226), .B(N2308), .S(net723969), .Q(n3519) );
  NAND24 U4008 ( .A(n3205), .B(n3206), .Q(net716181) );
  INV6 U4009 ( .A(n2865), .Q(n3846) );
  INV1 U4010 ( .A(net712607), .Q(net723758) );
  XNR20 U4011 ( .A(net712952), .B(net715576), .Q(net712965) );
  NAND26 U4012 ( .A(net712939), .B(net712940), .Q(net712952) );
  CLKIN6 U4013 ( .A(net712945), .Q(net718373) );
  INV10 U4014 ( .A(n3727), .Q(n3737) );
  INV0 U4015 ( .A(n3297), .Q(n3207) );
  CLKIN12 U4016 ( .A(n3858), .Q(n3872) );
  INV12 U4017 ( .A(n3673), .Q(n3722) );
  NAND24 U4018 ( .A(n3256), .B(net715678), .Q(net712950) );
  XNR22 U4019 ( .A(net712993), .B(n3629), .Q(n3256) );
  XOR22 U4020 ( .A(n3658), .B(net725513), .Q(n3659) );
  AOI212 U4021 ( .A(n3291), .B(net725513), .C(n3972), .Q(n3983) );
  NAND28 U4022 ( .A(n3224), .B(n3225), .Q(net724837) );
  NAND24 U4023 ( .A(net712888), .B(net715450), .Q(n3666) );
  NAND22 U4024 ( .A(n3429), .B(net712166), .Q(net725472) );
  INV3 U4025 ( .A(net725472), .Q(net725473) );
  NAND28 U4026 ( .A(n3210), .B(net725460), .Q(n3212) );
  NAND28 U4027 ( .A(n3211), .B(n3212), .Q(net721166) );
  INV2 U4028 ( .A(net712871), .Q(net725460) );
  INV6 U4029 ( .A(n3650), .Q(n3210) );
  INV1 U4030 ( .A(net720041), .Q(net725453) );
  INV0 U4031 ( .A(net715768), .Q(net720041) );
  NAND24 U4032 ( .A(net720042), .B(net725448), .Q(n3216) );
  INV1 U4033 ( .A(net723912), .Q(net725448) );
  NAND28 U4034 ( .A(n3218), .B(n4119), .Q(n4282) );
  INV1 U4035 ( .A(n3554), .Q(n4120) );
  NAND22 U4036 ( .A(n3620), .B(n3619), .Q(n3220) );
  NAND28 U4037 ( .A(n3623), .B(n3219), .Q(n3221) );
  NOR23 U4038 ( .A(n3223), .B(n3707), .Q(n3710) );
  INV1 U4039 ( .A(net723472), .Q(net725419) );
  NAND33 U4040 ( .A(net712877), .B(net719152), .C(n3656), .Q(n3677) );
  INV12 U4041 ( .A(net713101), .Q(net713073) );
  NAND26 U4042 ( .A(n3617), .B(net713041), .Q(n3621) );
  AOI311 U4043 ( .A(n3627), .B(net713005), .C(n3626), .D(n3625), .Q(n3628) );
  BUF15 U4044 ( .A(n4281), .Q(n3544) );
  NAND24 U4045 ( .A(N2475), .B(net718129), .Q(n4098) );
  NAND21 U4046 ( .A(net722521), .B(N2966), .Q(n4210) );
  CLKIN6 U4047 ( .A(net717664), .Q(net719771) );
  NAND22 U4048 ( .A(net718162), .B(N2666), .Q(n4121) );
  INV6 U4049 ( .A(n4133), .Q(n4103) );
  NAND24 U4050 ( .A(N2559), .B(net715360), .Q(n4133) );
  NAND23 U4051 ( .A(n3373), .B(n3766), .Q(n3753) );
  INV6 U4052 ( .A(n4053), .Q(n4250) );
  MUX24 U4053 ( .A(N2101), .B(net723498), .S(net712079), .Q(n3227) );
  BUF15 U4054 ( .A(net718011), .Q(net715717) );
  NAND26 U4055 ( .A(n3457), .B(n3456), .Q(net712646) );
  INV6 U4056 ( .A(net713181), .Q(net716401) );
  NAND32 U4057 ( .A(net723883), .B(net715576), .C(n2924), .Q(n3387) );
  INV0 U4058 ( .A(net715480), .Q(net719727) );
  BUF2 U4059 ( .A(net715674), .Q(net715825) );
  CLKIN8 U4060 ( .A(n4081), .Q(n4246) );
  MUX26 U4061 ( .A(N2116), .B(N1987), .S(n3577), .Q(n3226) );
  INV3 U4062 ( .A(net712513), .Q(net724864) );
  MUX26 U4063 ( .A(N2115), .B(N1986), .S(n3577), .Q(n3228) );
  MUX24 U4064 ( .A(n3228), .B(N2307), .S(net723969), .Q(n3229) );
  INV0 U4065 ( .A(net721373), .Q(net721134) );
  INV3 U4066 ( .A(arg[26]), .Q(net713170) );
  INV3 U4067 ( .A(n3424), .Q(n3425) );
  MUX26 U4068 ( .A(N1907), .B(n3529), .S(n2959), .Q(n3230) );
  INV0 U4069 ( .A(net712196), .Q(net723498) );
  MUX26 U4070 ( .A(N2104), .B(net721406), .S(n3578), .Q(n3231) );
  INV3 U4071 ( .A(n3940), .Q(n3415) );
  CLKIN6 U4072 ( .A(N1784), .Q(net716389) );
  INV3 U4073 ( .A(net723890), .Q(net712475) );
  INV1 U4074 ( .A(n3309), .Q(n3684) );
  XNR21 U4075 ( .A(net720185), .B(n3641), .Q(n3309) );
  INV3 U4076 ( .A(n3684), .Q(n3366) );
  INV3 U4077 ( .A(net724125), .Q(net712931) );
  CLKIN1 U4078 ( .A(net712957), .Q(net724125) );
  MUX22 U4079 ( .A(n4299), .B(N2277), .S(net715725), .Q(n3232) );
  NAND24 U4080 ( .A(net712793), .B(net718624), .Q(n3450) );
  INV6 U4081 ( .A(n3837), .Q(n3826) );
  BUF2 U4082 ( .A(net723541), .Q(net725181) );
  NAND26 U4083 ( .A(net712696), .B(net715769), .Q(net712559) );
  BUF2 U4084 ( .A(n3738), .Q(n3233) );
  NOR33 U4085 ( .A(n3804), .B(net715576), .C(net712493), .Q(n3805) );
  NAND24 U4086 ( .A(n3387), .B(n2944), .Q(n3718) );
  MUX26 U4087 ( .A(n3524), .B(N2305), .S(net715717), .Q(n3262) );
  NAND22 U4088 ( .A(net715753), .B(N2860), .Q(n4200) );
  NAND21 U4089 ( .A(N2878), .B(net722433), .Q(n4168) );
  CLKIN6 U4090 ( .A(n3875), .Q(n3730) );
  NAND24 U4091 ( .A(net712803), .B(net712793), .Q(n3685) );
  NAND24 U4092 ( .A(net712730), .B(net712729), .Q(n3393) );
  INV3 U4093 ( .A(net715788), .Q(net725117) );
  INV6 U4094 ( .A(net713148), .Q(net713138) );
  CLKIN3 U4095 ( .A(net713100), .Q(net713097) );
  INV2 U4096 ( .A(net713099), .Q(net713098) );
  NAND22 U4097 ( .A(n3348), .B(n3349), .Q(N2540) );
  AOI212 U4098 ( .A(net719298), .B(net723292), .C(n3553), .Q(n3235) );
  OAI212 U4099 ( .A(net713067), .B(net713068), .C(n3432), .Q(net713066) );
  AOI2112 U4100 ( .A(net726165), .B(n3531), .C(n4020), .D(n4019), .Q(net712168) );
  CLKIN6 U4101 ( .A(n4087), .Q(N2550) );
  IMUX21 U4102 ( .A(n2863), .B(N2491), .S(net717907), .Q(n4082) );
  NOR24 U4103 ( .A(net724923), .B(net719237), .Q(n3237) );
  NAND26 U4104 ( .A(n3317), .B(arg[17]), .Q(n3319) );
  BUF2 U4105 ( .A(n3239), .Q(n3238) );
  NAND33 U4106 ( .A(n3372), .B(net724188), .C(net724863), .Q(n3373) );
  CLKIN6 U4107 ( .A(n3459), .Q(n3460) );
  BUF15 U4108 ( .A(N2548), .Q(n3555) );
  NAND20 U4109 ( .A(n3801), .B(net715572), .Q(n3803) );
  MUX24 U4110 ( .A(N2094), .B(n3531), .S(net712079), .Q(n3239) );
  BUF2 U4111 ( .A(n3528), .Q(n3240) );
  NAND21 U4112 ( .A(n3871), .B(n3297), .Q(n3859) );
  BUF2 U4113 ( .A(N2553), .Q(n3241) );
  INV6 U4114 ( .A(n3760), .Q(n3761) );
  NAND22 U4115 ( .A(n3695), .B(net712712), .Q(n3318) );
  NAND24 U4116 ( .A(net724795), .B(net715788), .Q(n3943) );
  NAND30 U4117 ( .A(net712877), .B(net719152), .C(n3656), .Q(n3243) );
  OAI222 U4118 ( .A(net723917), .B(n3802), .C(net712496), .D(n3803), .Q(n3806)
         );
  INV2 U4119 ( .A(n3565), .Q(n3567) );
  INV2 U4120 ( .A(n3782), .Q(n3778) );
  XNR22 U4121 ( .A(net715775), .B(n3568), .Q(n3868) );
  CLKIN6 U4122 ( .A(n3911), .Q(n3568) );
  NAND28 U4123 ( .A(n3318), .B(n3319), .Q(net712710) );
  NAND28 U4124 ( .A(n3455), .B(net718580), .Q(n3457) );
  NAND22 U4125 ( .A(net717664), .B(N2669), .Q(n4115) );
  OAI222 U4126 ( .A(N2688), .B(n4103), .C(net722561), .D(n4103), .Q(n4104) );
  NAND28 U4127 ( .A(net716402), .B(net724167), .Q(net710022) );
  XOR20 U4128 ( .A(net721834), .B(n3233), .Q(n3244) );
  BUF2 U4129 ( .A(net712567), .Q(net724758) );
  NAND28 U4130 ( .A(net715480), .B(net712917), .Q(n3635) );
  XNR22 U4131 ( .A(net715769), .B(n3639), .Q(n3640) );
  OAI2112 U4132 ( .A(n3595), .B(n3594), .C(net713166), .D(net715768), .Q(n3245) );
  OAI311 U4133 ( .A(net719616), .B(arg[31]), .C(net720121), .D(net713184), .Q(
        n3595) );
  NAND22 U4134 ( .A(N2673), .B(net717664), .Q(n4111) );
  NAND34 U4135 ( .A(n3236), .B(n3389), .C(n3885), .Q(n3248) );
  NAND32 U4136 ( .A(n3236), .B(n3389), .C(n3885), .Q(n3890) );
  CLKIN3 U4137 ( .A(net719771), .Q(net724671) );
  CLKIN2 U4138 ( .A(net724795), .Q(net723444) );
  INV12 U4139 ( .A(net712214), .Q(N1781) );
  CLKIN1 U4140 ( .A(n3690), .Q(n3295) );
  CLKIN6 U4141 ( .A(n3729), .Q(n3250) );
  INV0 U4142 ( .A(n3729), .Q(n3877) );
  XNR22 U4143 ( .A(n3736), .B(net721373), .Q(n3253) );
  NAND26 U4144 ( .A(n3971), .B(n3392), .Q(n3986) );
  INV6 U4145 ( .A(n3564), .Q(n3251) );
  CLKIN6 U4146 ( .A(n3964), .Q(n3564) );
  XNR22 U4147 ( .A(net724508), .B(n3844), .Q(net712434) );
  INV3 U4148 ( .A(net712677), .Q(net721162) );
  INV2 U4149 ( .A(n3772), .Q(n3252) );
  INV1 U4150 ( .A(n3771), .Q(n3772) );
  NAND21 U4151 ( .A(net712612), .B(net715712), .Q(n3771) );
  XOR22 U4152 ( .A(n3789), .B(net712475), .Q(n3274) );
  NOR42 U4153 ( .A(n3969), .B(n3251), .C(n3942), .D(n3290), .Q(n3953) );
  CLKIN4 U4154 ( .A(n3773), .Q(n3254) );
  INV6 U4155 ( .A(n3254), .Q(n3255) );
  CLKIN0 U4156 ( .A(net712145), .Q(net721406) );
  IMUX23 U4157 ( .A(n3328), .B(net723106), .S(n3578), .Q(n3305) );
  INV12 U4158 ( .A(n4012), .Q(N1779) );
  CLKIN0 U4159 ( .A(n3801), .Q(n3257) );
  CLKIN6 U4160 ( .A(n3815), .Q(n3801) );
  BUF2 U4161 ( .A(net716181), .Q(net723959) );
  MUX26 U4162 ( .A(n4237), .B(N2474), .S(net717907), .Q(n3258) );
  INV0 U4163 ( .A(n4243), .Q(n3259) );
  NAND22 U4164 ( .A(n3270), .B(n3949), .Q(n3383) );
  BUF2 U4165 ( .A(n4222), .Q(n3260) );
  MUX24 U4166 ( .A(N2297), .B(n3513), .S(net719234), .Q(n3261) );
  BUF2 U4167 ( .A(n2872), .Q(net724508) );
  INV3 U4168 ( .A(n4249), .Q(n3263) );
  MUX26 U4169 ( .A(n3337), .B(N2100), .S(n3575), .Q(n3264) );
  INV6 U4170 ( .A(net712655), .Q(net712654) );
  NAND24 U4171 ( .A(n3265), .B(net715544), .Q(n3930) );
  XOR22 U4172 ( .A(net712536), .B(n3790), .Q(n3265) );
  INV6 U4173 ( .A(n3767), .Q(n3774) );
  NAND24 U4174 ( .A(net718090), .B(n2903), .Q(n4070) );
  INV6 U4175 ( .A(N2293), .Q(n4060) );
  INV0 U4176 ( .A(n2862), .Q(n3266) );
  INV0 U4177 ( .A(n4223), .Q(n4197) );
  XNR22 U4178 ( .A(n3738), .B(net721834), .Q(n3267) );
  INV6 U4179 ( .A(n3743), .Q(n3427) );
  NAND24 U4180 ( .A(net712732), .B(net712760), .Q(n3695) );
  INV4 U4181 ( .A(n3842), .Q(n3493) );
  NAND26 U4182 ( .A(n3493), .B(net718362), .Q(n3495) );
  OAI212 U4183 ( .A(net720567), .B(n3569), .C(n3910), .Q(n3912) );
  NOR33 U4184 ( .A(n3425), .B(n3507), .C(net716172), .Q(n3910) );
  INV3 U4185 ( .A(n3764), .Q(n3747) );
  NAND26 U4186 ( .A(n3359), .B(n3358), .Q(n3361) );
  INV3 U4187 ( .A(n3900), .Q(n3359) );
  INV1 U4188 ( .A(n3272), .Q(n3270) );
  OAI312 U4189 ( .A(net712582), .B(n3765), .C(net720253), .D(n3756), .Q(n3760)
         );
  NAND22 U4190 ( .A(n3914), .B(net715700), .Q(n4011) );
  BUF2 U4191 ( .A(N1785), .Q(n3396) );
  NAND23 U4192 ( .A(n3900), .B(n3507), .Q(n3360) );
  INV6 U4193 ( .A(N1793), .Q(n3284) );
  NOR42 U4194 ( .A(n3970), .B(n3972), .C(n3951), .D(n3199), .Q(n3952) );
  OAI222 U4195 ( .A(n3846), .B(n3847), .C(n3543), .D(n3845), .Q(n3851) );
  XOR22 U4196 ( .A(n3811), .B(net725181), .Q(n3272) );
  OAI222 U4197 ( .A(net723273), .B(net712454), .C(arg[14]), .D(n3925), .Q(
        n3941) );
  XNR22 U4198 ( .A(n3990), .B(n4001), .Q(n3273) );
  OAI312 U4199 ( .A(arg[27]), .B(n3601), .C(net713090), .D(n3600), .Q(n3602)
         );
  OAI212 U4200 ( .A(net712369), .B(n3897), .C(n3896), .Q(n3944) );
  NAND26 U4201 ( .A(net722414), .B(net716402), .Q(net713129) );
  INV1 U4202 ( .A(net712918), .Q(net723674) );
  OAI212 U4203 ( .A(net721379), .B(n3728), .C(net715540), .Q(n3729) );
  CLKIN0 U4204 ( .A(net712698), .Q(net723751) );
  BUF2 U4205 ( .A(net712573), .Q(net723881) );
  NAND28 U4206 ( .A(n4010), .B(n3284), .Q(n3917) );
  OAI222 U4207 ( .A(n3236), .B(n3839), .C(net725513), .D(n2864), .Q(n3841) );
  OAI212 U4208 ( .A(net712369), .B(n3897), .C(n3896), .Q(n3276) );
  NAND33 U4209 ( .A(arg[28]), .B(net719607), .C(arg[30]), .Q(net723781) );
  NAND22 U4210 ( .A(n4233), .B(net719447), .Q(net711940) );
  INV3 U4211 ( .A(n3800), .Q(n3474) );
  INV6 U4212 ( .A(net722413), .Q(net724167) );
  INV10 U4213 ( .A(n3546), .Q(n4208) );
  NAND28 U4214 ( .A(n3622), .B(n3621), .Q(n3626) );
  NAND24 U4215 ( .A(net712903), .B(net715768), .Q(net713005) );
  NAND20 U4216 ( .A(n3812), .B(net715608), .Q(n3799) );
  OAI212 U4217 ( .A(net722561), .B(n3395), .C(n4105), .Q(n3277) );
  CLKIN3 U4218 ( .A(net713125), .Q(net713130) );
  BUF2 U4219 ( .A(net713011), .Q(net724119) );
  NAND24 U4220 ( .A(net715480), .B(n3626), .Q(n3412) );
  AOI212 U4221 ( .A(n2877), .B(n3426), .C(net712877), .Q(n3281) );
  INV4 U4222 ( .A(net712904), .Q(net713074) );
  CLKIN6 U4223 ( .A(net713162), .Q(net723251) );
  XNR22 U4224 ( .A(net715572), .B(n3853), .Q(n3854) );
  NOR22 U4225 ( .A(net712211), .B(n3931), .Q(n3933) );
  NOR23 U4226 ( .A(net712123), .B(net712124), .Q(n3283) );
  NAND21 U4227 ( .A(n3928), .B(n3929), .Q(n3945) );
  NOR23 U4228 ( .A(N1985), .B(N1978), .Q(net712125) );
  CLKIN6 U4229 ( .A(net713161), .Q(net722413) );
  AOI222 U4230 ( .A(n3950), .B(net715616), .C(n3830), .D(net715576), .Q(n3827)
         );
  XOR22 U4231 ( .A(net715576), .B(n3651), .Q(n3652) );
  IMUX20 U4232 ( .A(net715680), .B(n3286), .S(net722521), .Q(sqroot[13]) );
  NAND21 U4233 ( .A(n3309), .B(n3724), .Q(n3671) );
  INV2 U4234 ( .A(net712792), .Q(net721256) );
  XOR22 U4235 ( .A(net715788), .B(net712305), .Q(n3931) );
  CLKIN0 U4236 ( .A(n3380), .Q(n4114) );
  OAI222 U4237 ( .A(net725733), .B(n3338), .C(n3964), .D(n3963), .Q(n3965) );
  NAND21 U4238 ( .A(n3529), .B(net715544), .Q(n3963) );
  INV0 U4239 ( .A(n3261), .Q(n3287) );
  BUF2 U4240 ( .A(net712415), .Q(net723961) );
  OAI212 U4241 ( .A(n3311), .B(n2934), .C(n3869), .Q(n3870) );
  INV1 U4242 ( .A(n3569), .Q(n3311) );
  INV0 U4243 ( .A(n2924), .Q(n3288) );
  NAND26 U4244 ( .A(n3573), .B(n3985), .Q(n3989) );
  NAND26 U4245 ( .A(n3369), .B(net722174), .Q(n3371) );
  CLKIN6 U4246 ( .A(n3755), .Q(n3369) );
  IMUX24 U4247 ( .A(n3768), .B(n3769), .S(net723927), .Q(n3770) );
  INV6 U4248 ( .A(n3836), .Q(n3848) );
  INV0 U4249 ( .A(n4238), .Q(n3289) );
  CLKIN8 U4250 ( .A(n4039), .Q(N1971) );
  NAND28 U4251 ( .A(n3370), .B(n3371), .Q(n3785) );
  INV2 U4252 ( .A(N1783), .Q(n3291) );
  CLKIN0 U4253 ( .A(n3757), .Q(n3292) );
  XNR22 U4254 ( .A(net723891), .B(n3789), .Q(n3566) );
  CLKIN2 U4255 ( .A(n3992), .Q(n3293) );
  NAND22 U4256 ( .A(n3755), .B(net723751), .Q(n3370) );
  BUF2 U4257 ( .A(n3253), .Q(n3294) );
  XOR22 U4258 ( .A(n3693), .B(n3295), .Q(net723873) );
  NAND21 U4259 ( .A(net720329), .B(n3421), .Q(n3422) );
  INV3 U4260 ( .A(net719771), .Q(net723850) );
  CLKIN0 U4261 ( .A(n3550), .Q(n4195) );
  CLKIN0 U4262 ( .A(n3400), .Q(n4118) );
  CLKIN15 U4263 ( .A(net719327), .Q(net718128) );
  INV12 U4264 ( .A(n3694), .Q(n3690) );
  AOI211 U4265 ( .A(net723758), .B(net712596), .C(net712610), .Q(n3756) );
  INV4 U4266 ( .A(net712991), .Q(net712895) );
  NAND24 U4267 ( .A(n3852), .B(n3471), .Q(n3472) );
  INV2 U4268 ( .A(net712501), .Q(net718466) );
  NOR40 U4269 ( .A(n3905), .B(n3906), .C(net723637), .D(n3873), .Q(n3874) );
  NOR30 U4270 ( .A(n3906), .B(net723637), .C(n3905), .Q(n3907) );
  CLKIN3 U4271 ( .A(n3906), .Q(n3314) );
  INV2 U4272 ( .A(n3905), .Q(n3780) );
  NOR24 U4273 ( .A(net715576), .B(n3686), .Q(net712777) );
  INV3 U4274 ( .A(net712644), .Q(net712680) );
  NAND22 U4275 ( .A(net712991), .B(net719166), .Q(net719165) );
  CLKIN6 U4276 ( .A(net712752), .Q(net712753) );
  BUF2 U4277 ( .A(n3858), .Q(n3297) );
  XNR22 U4278 ( .A(net712782), .B(n3687), .Q(n3702) );
  NAND23 U4279 ( .A(n3761), .B(net725513), .Q(n3386) );
  NAND21 U4280 ( .A(net712415), .B(n3297), .Q(n3905) );
  NOR21 U4281 ( .A(net721242), .B(n3667), .Q(n3668) );
  INV1 U4282 ( .A(n3666), .Q(n3667) );
  INV3 U4283 ( .A(n3671), .Q(n3672) );
  NAND22 U4284 ( .A(N2556), .B(net715360), .Q(n4139) );
  NAND33 U4285 ( .A(n3737), .B(net715540), .C(n3726), .Q(n3875) );
  NOR41 U4286 ( .A(n3776), .B(n3732), .C(net721379), .D(n3731), .Q(n3726) );
  AOI312 U4287 ( .A(net712605), .B(net723768), .C(net712596), .D(n3749), .Q(
        n3750) );
  MUX24 U4288 ( .A(N2296), .B(n3231), .S(net719234), .Q(n3298) );
  BUF2 U4289 ( .A(n4292), .Q(n3299) );
  BUF2 U4290 ( .A(N2546), .Q(n3300) );
  CLKIN0 U4291 ( .A(n4240), .Q(n3301) );
  CLKIN0 U4292 ( .A(n3516), .Q(n3302) );
  INV3 U4293 ( .A(n3302), .Q(n3303) );
  BUF2 U4294 ( .A(N2544), .Q(n3304) );
  NAND22 U4295 ( .A(n3935), .B(n3415), .Q(n3416) );
  INV1 U4296 ( .A(n4210), .Q(sqroot[16]) );
  NOR24 U4297 ( .A(n3307), .B(net719237), .Q(n3306) );
  XNR22 U4298 ( .A(net715678), .B(n3638), .Q(n3633) );
  NAND24 U4299 ( .A(n3272), .B(net715608), .Q(n3849) );
  NAND24 U4300 ( .A(n3352), .B(n3353), .Q(net712483) );
  OAI222 U4301 ( .A(arg[18]), .B(n3691), .C(n2872), .D(n3690), .Q(net723555)
         );
  OAI210 U4302 ( .A(net712760), .B(net715542), .C(net712531), .Q(n3308) );
  AOI2112 U4303 ( .A(net712743), .B(n3701), .C(net723702), .D(net712744), .Q(
        n3704) );
  AOI212 U4304 ( .A(arg[27]), .B(arg[26]), .C(net713211), .Q(net723527) );
  NAND23 U4305 ( .A(n3587), .B(n3586), .Q(net713211) );
  AOI222 U4306 ( .A(net712983), .B(net712984), .C(net712985), .D(net716699), 
        .Q(net723514) );
  NAND21 U4307 ( .A(n3624), .B(net724119), .Q(net713001) );
  CLKIN0 U4308 ( .A(n2899), .Q(n3312) );
  AOI222 U4309 ( .A(net716699), .B(net715712), .C(net712914), .D(net718388), 
        .Q(n3637) );
  CLKIN0 U4310 ( .A(net712885), .Q(net712871) );
  MUX24 U4311 ( .A(N2299), .B(n4253), .S(net719234), .Q(n3440) );
  INV12 U4312 ( .A(net702066), .Q(net715542) );
  CLKIN0 U4313 ( .A(n3830), .Q(n3313) );
  INV6 U4314 ( .A(n3677), .Q(n3664) );
  NAND26 U4315 ( .A(n4073), .B(n4072), .Q(n4093) );
  NAND24 U4316 ( .A(net718011), .B(n4062), .Q(n4072) );
  NAND24 U4317 ( .A(n3340), .B(net718090), .Q(n4073) );
  NAND22 U4318 ( .A(n3245), .B(net713162), .Q(n3321) );
  INV3 U4319 ( .A(n3596), .Q(n3320) );
  IMUX23 U4320 ( .A(n3514), .B(N2302), .S(net715717), .Q(n4079) );
  INV10 U4321 ( .A(net720894), .Q(net722482) );
  NAND24 U4322 ( .A(n3316), .B(n3783), .Q(net712544) );
  INV3 U4323 ( .A(n3784), .Q(n3315) );
  INV2 U4324 ( .A(n3913), .Q(n3914) );
  NAND24 U4325 ( .A(n3321), .B(n3322), .Q(net713159) );
  NAND24 U4326 ( .A(n3431), .B(n3430), .Q(n3768) );
  BUF2 U4327 ( .A(n4239), .Q(n3323) );
  NAND24 U4328 ( .A(N2686), .B(net722561), .Q(n4137) );
  CLKIN1 U4329 ( .A(n3270), .Q(n3381) );
  INV0 U4330 ( .A(n3305), .Q(n3340) );
  BUF2 U4331 ( .A(n2925), .Q(n3324) );
  CLKIN6 U4332 ( .A(n3598), .Q(n3597) );
  INV2 U4333 ( .A(n3883), .Q(n3389) );
  INV6 U4334 ( .A(n4070), .Q(n4059) );
  NAND22 U4335 ( .A(n4140), .B(n4139), .Q(n4265) );
  BUF2 U4336 ( .A(n3203), .Q(n3325) );
  NAND23 U4337 ( .A(net718471), .B(n3473), .Q(net718473) );
  NAND23 U4338 ( .A(n3530), .B(net721041), .Q(n4158) );
  NAND23 U4339 ( .A(net724065), .B(net713058), .Q(n3620) );
  NAND22 U4340 ( .A(net717815), .B(net717816), .Q(n3583) );
  BUF2 U4341 ( .A(net712518), .Q(net720787) );
  NAND21 U4342 ( .A(net720274), .B(N2868), .Q(n4187) );
  NAND20 U4343 ( .A(net715540), .B(n3790), .Q(n3791) );
  NAND23 U4344 ( .A(n3830), .B(net715576), .Q(n3882) );
  CLKIN4 U4345 ( .A(net715745), .Q(net720986) );
  CLKIN6 U4346 ( .A(net713103), .Q(net721341) );
  INV3 U4347 ( .A(net718617), .Q(net720826) );
  NAND26 U4348 ( .A(n3598), .B(net713114), .Q(net713057) );
  CLKIN1 U4349 ( .A(net713061), .Q(net718617) );
  NAND24 U4350 ( .A(n3406), .B(net711884), .Q(res_3_) );
  INV6 U4351 ( .A(n3670), .Q(n3682) );
  INV1 U4352 ( .A(n3289), .Q(n3355) );
  CLKIN2 U4353 ( .A(n4241), .Q(n3357) );
  NAND23 U4354 ( .A(n3948), .B(net712286), .Q(n3949) );
  MUX24 U4355 ( .A(n3331), .B(n3332), .S(net712079), .Q(n3330) );
  IMUX23 U4356 ( .A(N1911), .B(N1782), .S(n2959), .Q(net712114) );
  NAND28 U4357 ( .A(n3335), .B(n3336), .Q(n3529) );
  CLKIN6 U4358 ( .A(net721637), .Q(net722912) );
  BUF2 U4359 ( .A(net712316), .Q(net721637) );
  AOI312 U4360 ( .A(n3890), .B(net715480), .C(n2895), .D(n3888), .Q(n3895) );
  NAND20 U4361 ( .A(N1917), .B(net715402), .Q(n4047) );
  CLKIN0 U4362 ( .A(n3200), .Q(n3337) );
  AOI2112 U4363 ( .A(net721714), .B(net715816), .C(n3921), .D(n3962), .Q(n3924) );
  AOI312 U4364 ( .A(n3861), .B(net722889), .C(n3887), .D(n3860), .Q(n3862) );
  INV0 U4365 ( .A(net723419), .Q(net718580) );
  NAND24 U4366 ( .A(N1906), .B(net725944), .Q(n3342) );
  CLKIN8 U4367 ( .A(n4009), .Q(N1790) );
  MUX24 U4368 ( .A(N2112), .B(N1983), .S(n3577), .Q(n3339) );
  NAND28 U4369 ( .A(n3383), .B(n3384), .Q(N1782) );
  NAND26 U4370 ( .A(n3382), .B(n3381), .Q(n3384) );
  OAI212 U4371 ( .A(net715768), .B(net720042), .C(net726021), .Q(n3769) );
  IMUX22 U4372 ( .A(N2099), .B(n2898), .S(net712079), .Q(n4053) );
  AOI212 U4373 ( .A(n3892), .B(net715711), .C(net720318), .Q(n3897) );
  NAND28 U4374 ( .A(n3342), .B(n3343), .Q(net722738) );
  INV1 U4375 ( .A(n3978), .Q(n3898) );
  NAND28 U4376 ( .A(n3934), .B(n3462), .Q(net712214) );
  NAND23 U4377 ( .A(net712175), .B(net720783), .Q(n4023) );
  AOI222 U4378 ( .A(net722729), .B(net716101), .C(N1968), .D(net723637), .Q(
        n3344) );
  OAI212 U4379 ( .A(net715480), .B(n3889), .C(net712369), .Q(n3888) );
  CLKIN0 U4380 ( .A(n3265), .Q(n3419) );
  BUF2 U4381 ( .A(n3555), .Q(n3345) );
  INV0 U4382 ( .A(n4272), .Q(n4186) );
  NAND22 U4383 ( .A(net722422), .B(n4246), .Q(n3458) );
  IMUX22 U4384 ( .A(n3339), .B(N2304), .S(net722482), .Q(n4055) );
  CLKBU12 U4385 ( .A(N2627), .Q(net715739) );
  NAND22 U4386 ( .A(net717664), .B(N2664), .Q(n4122) );
  OAI212 U4387 ( .A(net719548), .B(n4175), .C(n4174), .Q(res_22_) );
  NAND23 U4388 ( .A(N2684), .B(net724671), .Q(n4142) );
  NAND22 U4389 ( .A(N2883), .B(net719548), .Q(n4162) );
  INV6 U4390 ( .A(net712700), .Q(net712789) );
  NAND28 U4391 ( .A(n3720), .B(n3719), .Q(n3727) );
  NOR41 U4392 ( .A(n3776), .B(n3732), .C(n3731), .D(n3727), .Q(n3728) );
  MUX21 U4393 ( .A(net726169), .B(N2956), .S(net711876), .Q(sqroot[6]) );
  NAND22 U4394 ( .A(n3721), .B(net721315), .Q(n3511) );
  OAI212 U4395 ( .A(net719548), .B(n4169), .C(n4168), .Q(res_25_) );
  INV6 U4396 ( .A(n4089), .Q(n4290) );
  CLKIN3 U4397 ( .A(N2627), .Q(net715362) );
  INV3 U4398 ( .A(N2243), .Q(net715326) );
  INV12 U4399 ( .A(n3547), .Q(n3548) );
  INV4 U4400 ( .A(n4182), .Q(n4183) );
  INV0 U4401 ( .A(n3345), .Q(n4108) );
  NAND24 U4402 ( .A(N2676), .B(net717664), .Q(n4109) );
  INV6 U4403 ( .A(N2557), .Q(n3346) );
  CLKIN12 U4404 ( .A(n3346), .Q(n3347) );
  INV6 U4405 ( .A(n4109), .Q(n3557) );
  NAND21 U4406 ( .A(N2873), .B(net719548), .Q(n4178) );
  NAND21 U4407 ( .A(N2882), .B(net719548), .Q(n4164) );
  NAND28 U4408 ( .A(n3348), .B(n3349), .Q(n3350) );
  NAND23 U4409 ( .A(N2682), .B(net719772), .Q(n4145) );
  NAND22 U4410 ( .A(net723435), .B(n3351), .Q(n3352) );
  NAND22 U4411 ( .A(n3798), .B(net715788), .Q(n3353) );
  INV3 U4412 ( .A(n3798), .Q(n3351) );
  BUF15 U4413 ( .A(n4286), .Q(n3546) );
  CLKIN0 U4414 ( .A(n3304), .Q(n4112) );
  BUF15 U4415 ( .A(N2627), .Q(net717664) );
  MUX21 U4416 ( .A(n4258), .B(N2884), .S(net722433), .Q(res_31_) );
  NAND22 U4417 ( .A(n3500), .B(n3501), .Q(n3502) );
  NAND22 U4418 ( .A(N2879), .B(net719548), .Q(n4166) );
  NAND22 U4419 ( .A(N2482), .B(net718129), .Q(net712018) );
  CLKIN6 U4420 ( .A(n4016), .Q(N1978) );
  INV2 U4421 ( .A(n3439), .Q(n4188) );
  NAND26 U4422 ( .A(net722422), .B(n3355), .Q(n3356) );
  NAND28 U4423 ( .A(n3356), .B(n4098), .Q(N2538) );
  NAND22 U4424 ( .A(N2495), .B(net718226), .Q(n3453) );
  CLKIN2 U4425 ( .A(n3306), .Q(n3417) );
  OAI212 U4426 ( .A(net718226), .B(n3287), .C(n4085), .Q(N2552) );
  IMUX24 U4427 ( .A(net721443), .B(n3961), .S(net715416), .Q(n3397) );
  NAND21 U4428 ( .A(N2498), .B(net719306), .Q(n4074) );
  CLKIN1 U4429 ( .A(net724837), .Q(net718495) );
  INV2 U4430 ( .A(n3507), .Q(n3358) );
  NAND22 U4431 ( .A(n3660), .B(net723674), .Q(n3363) );
  NAND28 U4432 ( .A(n3363), .B(n3364), .Q(net712733) );
  CLKIN3 U4433 ( .A(net723674), .Q(net722234) );
  AOI2112 U4434 ( .A(net722222), .B(n3639), .C(net722223), .D(net715510), .Q(
        n3365) );
  INV12 U4435 ( .A(net712885), .Q(net712917) );
  INV6 U4436 ( .A(n3393), .Q(n3394) );
  AOI311 U4437 ( .A(n3308), .B(net712505), .C(net712512), .D(net712507), .Q(
        n3800) );
  BUF2 U4438 ( .A(n3757), .Q(n3368) );
  INV3 U4439 ( .A(n3752), .Q(n3372) );
  NAND24 U4440 ( .A(n2924), .B(n3374), .Q(n3376) );
  INV6 U4441 ( .A(n3751), .Q(n3766) );
  NAND28 U4442 ( .A(n3762), .B(net725513), .Q(net712605) );
  OAI222 U4443 ( .A(arg[18]), .B(n3691), .C(net715705), .D(n3690), .Q(n3701)
         );
  INV3 U4444 ( .A(n3653), .Q(n3654) );
  NAND26 U4445 ( .A(n3480), .B(net718432), .Q(n3482) );
  NAND20 U4446 ( .A(N1924), .B(net715761), .Q(n4043) );
  NAND24 U4447 ( .A(net712700), .B(net715788), .Q(net712743) );
  BUF2 U4448 ( .A(n4288), .Q(n3379) );
  BUF2 U4449 ( .A(n3541), .Q(n3380) );
  CLKIN6 U4450 ( .A(n3949), .Q(n3382) );
  OAI212 U4451 ( .A(net712680), .B(n3718), .C(n3717), .Q(n3719) );
  OAI222 U4452 ( .A(arg[18]), .B(n3691), .C(n2872), .D(n3690), .Q(net721808)
         );
  IMUX22 U4453 ( .A(n3867), .B(n3868), .S(n3399), .Q(n3869) );
  NAND21 U4454 ( .A(net712475), .B(net712139), .Q(n3817) );
  CLKIN6 U4455 ( .A(n3845), .Q(n3388) );
  OAI212 U4456 ( .A(net715825), .B(n3761), .C(net721638), .Q(n3763) );
  XNR21 U4457 ( .A(n3877), .B(n3874), .Q(n3996) );
  NAND28 U4458 ( .A(net712414), .B(net715825), .Q(n3887) );
  XNR22 U4459 ( .A(n3912), .B(n3390), .Q(n3526) );
  CLKIN6 U4460 ( .A(n4035), .Q(N1985) );
  NAND28 U4461 ( .A(n3510), .B(net717806), .Q(n3512) );
  NOR24 U4462 ( .A(n3391), .B(n3715), .Q(n3720) );
  NAND26 U4463 ( .A(net720274), .B(N2864), .Q(n4194) );
  INV4 U4464 ( .A(n4184), .Q(n4229) );
  INV0 U4465 ( .A(n3249), .Q(n4153) );
  IMUX20 U4466 ( .A(n4298), .B(N2278), .S(net723969), .Q(n4125) );
  INV0 U4467 ( .A(N2549), .Q(n3395) );
  NAND28 U4468 ( .A(n3414), .B(net720697), .Q(net720700) );
  XOR22 U4469 ( .A(n3753), .B(net719727), .Q(n3754) );
  NAND22 U4470 ( .A(N2680), .B(net722561), .Q(n4149) );
  INV4 U4471 ( .A(n3959), .Q(n3972) );
  NOR33 U4472 ( .A(n3970), .B(n3969), .C(n3968), .Q(n3971) );
  INV6 U4473 ( .A(n3616), .Q(n3622) );
  NAND28 U4474 ( .A(n3494), .B(n3495), .Q(N1784) );
  NAND21 U4475 ( .A(n3427), .B(net724008), .Q(net720124) );
  NAND26 U4476 ( .A(n3444), .B(n3445), .Q(net712905) );
  NOR22 U4477 ( .A(net712211), .B(n3936), .Q(n3937) );
  NAND21 U4478 ( .A(n3241), .B(net719447), .Q(n4146) );
  INV0 U4479 ( .A(N1777), .Q(net719965) );
  NAND22 U4480 ( .A(net718162), .B(n4126), .Q(n4160) );
  INV12 U4481 ( .A(arg[30]), .Q(net720121) );
  INV12 U4482 ( .A(arg[30]), .Q(net717815) );
  INV12 U4483 ( .A(arg[30]), .Q(net719952) );
  BUF15 U4484 ( .A(n4273), .Q(n3552) );
  INV3 U4485 ( .A(n4021), .Q(n4022) );
  NAND26 U4486 ( .A(n3398), .B(n3624), .Q(net713101) );
  INV2 U4487 ( .A(n3775), .Q(n3731) );
  AOI312 U4488 ( .A(n3426), .B(n3442), .C(n3656), .D(n3655), .Q(n3658) );
  CLKIN3 U4489 ( .A(net713097), .Q(net721349) );
  NAND33 U4490 ( .A(net720951), .B(net721340), .C(net721341), .Q(n3398) );
  INV2 U4491 ( .A(net715767), .Q(net721340) );
  NAND24 U4492 ( .A(net713104), .B(n3600), .Q(n3624) );
  CLKIN6 U4493 ( .A(n3829), .Q(n3498) );
  NOR42 U4494 ( .A(n3714), .B(n3222), .C(net725513), .D(net712721), .Q(n3709)
         );
  XOR22 U4495 ( .A(net715570), .B(n3698), .Q(n3699) );
  XOR22 U4496 ( .A(n3648), .B(net715478), .Q(n3649) );
  XNR22 U4497 ( .A(net715450), .B(n3427), .Q(n3742) );
  BUF2 U4498 ( .A(net712344), .Q(net721293) );
  NAND24 U4499 ( .A(n4147), .B(n4148), .Q(n4269) );
  NAND24 U4500 ( .A(n3458), .B(n4080), .Q(N2556) );
  INV3 U4501 ( .A(n4104), .Q(n4231) );
  BUF15 U4502 ( .A(net715346), .Q(net717907) );
  IMUX21 U4503 ( .A(n4248), .B(N2496), .S(net717907), .Q(n4077) );
  NAND22 U4504 ( .A(net718128), .B(N2478), .Q(n4096) );
  NOR24 U4505 ( .A(n4064), .B(n4063), .Q(n4242) );
  OAI221 U4506 ( .A(net715769), .B(net712903), .C(net713008), .D(net713009), 
        .Q(n3625) );
  OAI222 U4507 ( .A(n3401), .B(net712855), .C(net715572), .D(n3654), .Q(n3655)
         );
  NAND24 U4508 ( .A(n3451), .B(net712997), .Q(n3629) );
  CLKIN0 U4509 ( .A(net712810), .Q(net721077) );
  INV2 U4510 ( .A(net721077), .Q(net721078) );
  NAND24 U4511 ( .A(n3402), .B(net712931), .Q(n3403) );
  NAND28 U4512 ( .A(n3403), .B(n3404), .Q(net712885) );
  CLKIN0 U4513 ( .A(net712821), .Q(net721083) );
  NAND21 U4514 ( .A(N1915), .B(net725944), .Q(n4016) );
  NAND28 U4515 ( .A(net713055), .B(net713153), .Q(net713090) );
  BUF15 U4516 ( .A(net715376), .Q(net715754) );
  BUF12 U4517 ( .A(net715376), .Q(net715745) );
  BUF15 U4518 ( .A(net715376), .Q(net715746) );
  BUF2 U4519 ( .A(net712895), .Q(net721024) );
  XNR22 U4520 ( .A(net720693), .B(net721548), .Q(net721014) );
  NAND20 U4521 ( .A(net715362), .B(n3347), .Q(n4138) );
  NAND24 U4522 ( .A(net720986), .B(n3405), .Q(n3406) );
  NAND24 U4523 ( .A(n3486), .B(n3408), .Q(n3487) );
  INV6 U4524 ( .A(n3407), .Q(n3408) );
  NOR24 U4525 ( .A(n3409), .B(n3034), .Q(n3638) );
  CLKIN3 U4526 ( .A(n3638), .Q(n3486) );
  NAND28 U4527 ( .A(net713155), .B(n3597), .Q(net713058) );
  NAND26 U4528 ( .A(net713189), .B(net713171), .Q(n3591) );
  OAI212 U4529 ( .A(net715480), .B(net713078), .C(n3608), .Q(n3609) );
  NAND20 U4530 ( .A(n3779), .B(n3778), .Q(n3873) );
  AOI212 U4531 ( .A(n3697), .B(n2946), .C(net712751), .Q(n3698) );
  NAND28 U4532 ( .A(net718604), .B(net718343), .Q(n3497) );
  NAND24 U4533 ( .A(N2866), .B(net715746), .Q(n4191) );
  NAND22 U4534 ( .A(N2489), .B(net725641), .Q(n4085) );
  IMUX22 U4535 ( .A(n3379), .B(N2487), .S(net723620), .Q(n4087) );
  NAND24 U4536 ( .A(N2687), .B(net719772), .Q(n4135) );
  NOR33 U4537 ( .A(net712651), .B(net715542), .C(n3777), .Q(n3736) );
  NAND28 U4538 ( .A(n3481), .B(n3482), .Q(n3815) );
  CLKIN0 U4539 ( .A(net712503), .Q(net712502) );
  AOI312 U4540 ( .A(n3818), .B(n3817), .C(net715816), .D(n3816), .Q(n3823) );
  INV0 U4541 ( .A(net715480), .Q(net720727) );
  NAND24 U4542 ( .A(net712688), .B(net723883), .Q(net712775) );
  NAND26 U4543 ( .A(n3632), .B(net715576), .Q(net712938) );
  NAND22 U4544 ( .A(n3628), .B(net724738), .Q(net713002) );
  NAND22 U4545 ( .A(n3299), .B(net718090), .Q(n3508) );
  MUX24 U4546 ( .A(n3552), .B(N2869), .S(net715754), .Q(res_16_) );
  NAND28 U4547 ( .A(n3435), .B(n4194), .Q(res_11_) );
  NAND22 U4548 ( .A(n3901), .B(n2934), .Q(n3997) );
  INV3 U4549 ( .A(n4048), .Q(N1976) );
  MUX22 U4550 ( .A(N1921), .B(n3192), .S(net715406), .Q(n3520) );
  NOR22 U4551 ( .A(N1921), .B(N1918), .Q(n4025) );
  OAI212 U4552 ( .A(n3852), .B(n3851), .C(n3850), .Q(n3853) );
  NAND28 U4553 ( .A(n3939), .B(n3416), .Q(n4012) );
  BUF15 U4554 ( .A(n3941), .Q(n3543) );
  INV3 U4555 ( .A(n3882), .Q(n3861) );
  INV3 U4556 ( .A(n3848), .Q(n3471) );
  INV6 U4557 ( .A(n3556), .Q(n4274) );
  CLKBU12 U4558 ( .A(net712079), .Q(net715687) );
  CLKIN6 U4559 ( .A(n4095), .Q(n3418) );
  INV3 U4560 ( .A(n4095), .Q(n4241) );
  CLKIN0 U4561 ( .A(net721293), .Q(net720570) );
  BUF2 U4562 ( .A(net712341), .Q(net720567) );
  INV6 U4563 ( .A(n3967), .Q(n3964) );
  INV6 U4564 ( .A(n4071), .Q(n4289) );
  NAND22 U4565 ( .A(N2494), .B(net718226), .Q(n4078) );
  AOI222 U4566 ( .A(n3895), .B(n3894), .C(net712374), .D(n3893), .Q(n3896) );
  NAND22 U4567 ( .A(n3842), .B(net712414), .Q(n3494) );
  NAND23 U4568 ( .A(n3974), .B(net715572), .Q(n3959) );
  NAND22 U4569 ( .A(N2685), .B(net724671), .Q(n4140) );
  OAI212 U4570 ( .A(n2872), .B(n3484), .C(net706857), .Q(n3795) );
  AOI222 U4571 ( .A(n3442), .B(n3675), .C(n3279), .D(net712815), .Q(n3676) );
  NOR22 U4572 ( .A(net720401), .B(n3280), .Q(net720403) );
  INV3 U4573 ( .A(arg[28]), .Q(net720401) );
  XNR22 U4574 ( .A(arg[26]), .B(net710022), .Q(n3604) );
  CLKIN6 U4575 ( .A(n3976), .Q(n3969) );
  NAND24 U4576 ( .A(n4025), .B(n4024), .Q(n4029) );
  CLKBU15 U4577 ( .A(n4054), .Q(n3577) );
  IMUX24 U4578 ( .A(n3938), .B(n3937), .S(n3420), .Q(n3939) );
  NAND22 U4579 ( .A(N2865), .B(net715746), .Q(n4192) );
  NAND22 U4580 ( .A(net719964), .B(n3260), .Q(n4182) );
  NAND22 U4581 ( .A(n3422), .B(n4172), .Q(res_23_) );
  INV3 U4582 ( .A(n4173), .Q(n3421) );
  INV0 U4583 ( .A(n4215), .Q(n4173) );
  OAI212 U4584 ( .A(net721268), .B(n3266), .C(n4121), .Q(n3423) );
  INV6 U4585 ( .A(net712202), .Q(N1964) );
  NAND22 U4586 ( .A(net712286), .B(n3854), .Q(n3855) );
  NOR23 U4587 ( .A(n3232), .B(net715739), .Q(n3438) );
  BUF15 U4588 ( .A(net715374), .Q(net720274) );
  NOR20 U4589 ( .A(net712344), .B(net712216), .Q(n3424) );
  CLKBU8 U4590 ( .A(n3515), .Q(n3507) );
  XNR22 U4591 ( .A(n2874), .B(n3723), .Q(net712652) );
  NAND22 U4592 ( .A(n3367), .B(n3366), .Q(n3723) );
  INV3 U4593 ( .A(n3278), .Q(n3439) );
  INV3 U4594 ( .A(N1924), .Q(n4027) );
  INV6 U4595 ( .A(n3276), .Q(N1785) );
  NAND28 U4596 ( .A(n3733), .B(n3737), .Q(n3777) );
  NAND22 U4597 ( .A(N2683), .B(net719772), .Q(n4143) );
  INV6 U4598 ( .A(n3721), .Q(n3510) );
  NAND24 U4599 ( .A(net712478), .B(net712521), .Q(n3814) );
  OAI312 U4600 ( .A(net715678), .B(net715710), .C(n3607), .D(n3606), .Q(n3608)
         );
  BUF2 U4601 ( .A(net712905), .Q(net720185) );
  OAI222 U4602 ( .A(net719607), .B(net713189), .C(arg[29]), .D(arg[31]), .Q(
        n3582) );
  BUF15 U4603 ( .A(net715346), .Q(net719293) );
  NAND24 U4604 ( .A(n3944), .B(net715769), .Q(n3977) );
  NAND24 U4605 ( .A(n3746), .B(net712415), .Q(n3491) );
  INV0 U4606 ( .A(n4282), .Q(n4203) );
  NOR24 U4607 ( .A(N1979), .B(n4032), .Q(n4033) );
  INV3 U4608 ( .A(n3428), .Q(n3429) );
  OAI222 U4609 ( .A(net715719), .B(n4295), .C(N2281), .D(net720894), .Q(n4067)
         );
  IMUX24 U4610 ( .A(n4289), .B(N2486), .S(net719306), .Q(n4106) );
  NAND22 U4611 ( .A(net712568), .B(net715768), .Q(n3430) );
  NOR33 U4612 ( .A(n3714), .B(n3242), .C(n3713), .Q(n3715) );
  NAND24 U4613 ( .A(N2107), .B(n3576), .Q(n4051) );
  NOR42 U4614 ( .A(n3674), .B(net712816), .C(n3678), .D(n3401), .Q(n3675) );
  BUF2 U4615 ( .A(net720783), .Q(net715794) );
  INV2 U4616 ( .A(n4160), .Q(n4161) );
  NAND22 U4617 ( .A(n3696), .B(net712700), .Q(n3481) );
  INV3 U4618 ( .A(net719965), .Q(net719966) );
  INV15 U4619 ( .A(arg[30]), .Q(net719953) );
  NAND32 U4620 ( .A(net713189), .B(net719616), .C(net719952), .Q(n3587) );
  NOR33 U4621 ( .A(n3425), .B(n3507), .C(n3904), .Q(n3998) );
  INV3 U4622 ( .A(n3999), .Q(n4003) );
  XNR20 U4623 ( .A(n3661), .B(net715614), .Q(n3662) );
  INV1 U4624 ( .A(net724167), .Q(net713160) );
  BUF15 U4625 ( .A(N2543), .Q(n3541) );
  NAND22 U4626 ( .A(net715700), .B(arg[12]), .Q(n3920) );
  OAI222 U4627 ( .A(net715572), .B(n3974), .C(net715608), .D(net712214), .Q(
        n3975) );
  XNR22 U4628 ( .A(n4011), .B(net712216), .Q(n3916) );
  NAND24 U4629 ( .A(n3590), .B(net713194), .Q(net713151) );
  CLKIN12 U4630 ( .A(net712905), .Q(net713015) );
  OAI222 U4631 ( .A(n3758), .B(n3759), .C(n3410), .D(net712605), .Q(net712602)
         );
  AOI2112 U4632 ( .A(net715781), .B(net712145), .C(net715824), .D(net712146), 
        .Q(n4037) );
  OAI212 U4633 ( .A(net715769), .B(n3569), .C(net715700), .Q(n3867) );
  AOI212 U4634 ( .A(net712316), .B(net723637), .C(n3786), .Q(n3787) );
  NAND22 U4635 ( .A(net702066), .B(n3699), .Q(n3700) );
  AOI212 U4636 ( .A(net719606), .B(arg[30]), .C(arg[28]), .Q(n3593) );
  NAND34 U4637 ( .A(arg[28]), .B(net719607), .C(arg[30]), .Q(n3589) );
  NAND28 U4638 ( .A(net719606), .B(arg[30]), .Q(n3586) );
  INV2 U4639 ( .A(n3988), .Q(n3570) );
  CLKIN6 U4640 ( .A(n4208), .Q(n3437) );
  OAI212 U4641 ( .A(net715754), .B(n4181), .C(n4180), .Q(res_19_) );
  NAND22 U4642 ( .A(N2670), .B(net721268), .Q(n4156) );
  NAND21 U4643 ( .A(n3977), .B(N1784), .Q(n3979) );
  BUF2 U4644 ( .A(net712512), .Q(net719733) );
  XOR22 U4645 ( .A(net712782), .B(n3687), .Q(n3436) );
  CLKIN1 U4646 ( .A(net712842), .Q(net712782) );
  XOR22 U4647 ( .A(n3739), .B(net719727), .Q(n3705) );
  NAND20 U4648 ( .A(N1923), .B(net715759), .Q(n4044) );
  CLKIN6 U4649 ( .A(net713005), .Q(net713008) );
  NOR24 U4650 ( .A(net715542), .B(n3466), .Q(n3721) );
  INV6 U4651 ( .A(N2679), .Q(n4152) );
  NAND20 U4652 ( .A(net715348), .B(n4244), .Q(n4102) );
  NAND21 U4653 ( .A(net720274), .B(N2862), .Q(n4198) );
  INV6 U4654 ( .A(net712311), .Q(net712305) );
  INV15 U4655 ( .A(arg[28]), .Q(net719616) );
  INV15 U4656 ( .A(arg[31]), .Q(net719606) );
  INV15 U4657 ( .A(arg[31]), .Q(net719607) );
  INV15 U4658 ( .A(arg[31]), .Q(net719603) );
  INV4 U4659 ( .A(n3586), .Q(n3585) );
  INV15 U4660 ( .A(arg[31]), .Q(net713210) );
  NAND28 U4661 ( .A(arg[31]), .B(arg[30]), .Q(n3592) );
  MUX26 U4662 ( .A(N2110), .B(N1981), .S(net715687), .Q(n3514) );
  MUX26 U4663 ( .A(N2111), .B(n3525), .S(n3577), .Q(n3523) );
  MUX26 U4664 ( .A(N2113), .B(n3520), .S(n3577), .Q(n3524) );
  MUX24 U4665 ( .A(N2092), .B(n3533), .S(net712079), .Q(n4292) );
  CLKIN0 U4666 ( .A(n3259), .Q(n3473) );
  MUX24 U4667 ( .A(N1902), .B(arg[9]), .S(net715416), .Q(n3531) );
  OAI222 U4668 ( .A(net719548), .B(n4183), .C(N2871), .D(n4183), .Q(n4184) );
  BUF15 U4669 ( .A(net715745), .Q(net719548) );
  BUF15 U4670 ( .A(n4284), .Q(n3545) );
  INV1 U4671 ( .A(n4283), .Q(n4205) );
  MUX24 U4672 ( .A(n3521), .B(N2492), .S(n2867), .Q(n3517) );
  MUX26 U4673 ( .A(N2105), .B(N1976), .S(net715687), .Q(n3513) );
  NOR24 U4674 ( .A(n3438), .B(n4161), .Q(n4232) );
  OAI312 U4675 ( .A(n3905), .B(n3294), .C(n3906), .D(n3782), .Q(n3783) );
  NAND24 U4676 ( .A(n4145), .B(n4146), .Q(n4268) );
  OAI212 U4677 ( .A(n3748), .B(net712654), .C(n3771), .Q(n3735) );
  NOR31 U4678 ( .A(n3665), .B(n3279), .C(n3664), .Q(n3669) );
  INV15 U4679 ( .A(net718011), .Q(net718090) );
  NAND22 U4680 ( .A(net718162), .B(N2668), .Q(n4117) );
  MUX24 U4681 ( .A(n3502), .B(N2692), .S(net724671), .Q(n4258) );
  NAND22 U4682 ( .A(n3882), .B(net725513), .Q(n3839) );
  NAND22 U4683 ( .A(net712945), .B(arg[20]), .Q(n3489) );
  CLKIN12 U4684 ( .A(n4051), .Q(n4253) );
  OAI212 U4685 ( .A(net715360), .B(n4152), .C(n4151), .Q(n4271) );
  CLKBU15 U4686 ( .A(net715362), .Q(net719447) );
  XNR22 U4687 ( .A(n4236), .B(net718128), .Q(n4100) );
  INV6 U4688 ( .A(n4069), .Q(n4288) );
  CLKIN3 U4689 ( .A(n3438), .Q(n4159) );
  NAND23 U4690 ( .A(n4160), .B(n4159), .Q(n4209) );
  CLKIN6 U4691 ( .A(N2671), .Q(n4154) );
  NAND22 U4692 ( .A(n4155), .B(n4156), .Q(n4211) );
  INV3 U4693 ( .A(n4220), .Q(n4177) );
  NAND24 U4694 ( .A(n4146), .B(n4145), .Q(n4220) );
  NAND22 U4695 ( .A(N2677), .B(net715739), .Q(n4107) );
  NAND20 U4696 ( .A(N2500), .B(net718226), .Q(n3501) );
  NAND20 U4697 ( .A(n3519), .B(net718324), .Q(n3500) );
  INV0 U4698 ( .A(net721440), .Q(net711901) );
  NAND24 U4699 ( .A(N2108), .B(n3576), .Q(n4050) );
  BUF2 U4700 ( .A(n4250), .Q(n3441) );
  IMUX21 U4701 ( .A(n3262), .B(N2497), .S(net725641), .Q(n4076) );
  NAND22 U4702 ( .A(N2106), .B(n3576), .Q(n4052) );
  INV6 U4703 ( .A(n4090), .Q(n4243) );
  IMUX22 U4704 ( .A(n2902), .B(N2301), .S(net715719), .Q(n4081) );
  NAND21 U4705 ( .A(N2551), .B(net719447), .Q(n4150) );
  CLKIN6 U4706 ( .A(n4076), .Q(N2560) );
  CLKIN8 U4707 ( .A(n4050), .Q(n4254) );
  OAI212 U4708 ( .A(net715754), .B(n4197), .C(n4196), .Q(res_10_) );
  CLKIN6 U4709 ( .A(n4077), .Q(N2559) );
  CLKIN6 U4710 ( .A(n4079), .Q(n4247) );
  OAI212 U4711 ( .A(net715753), .B(n4201), .C(n4200), .Q(res_7_) );
  NAND22 U4712 ( .A(net715746), .B(N2858), .Q(n4204) );
  AOI212 U4713 ( .A(n3891), .B(net715712), .C(net712211), .Q(n3894) );
  OAI2112 U4714 ( .A(n3678), .B(n3243), .C(n3676), .D(net721078), .Q(n3679) );
  NOR42 U4715 ( .A(arg[30]), .B(arg[28]), .C(net713210), .D(arg[29]), .Q(n3580) );
  OAI221 U4716 ( .A(net721714), .B(net715816), .C(n3922), .D(net712323), .Q(
        n3923) );
  XNR22 U4717 ( .A(n4008), .B(n4007), .Q(n4009) );
  INV2 U4718 ( .A(n4217), .Q(n4175) );
  MUX24 U4719 ( .A(N2093), .B(N1964), .S(net712079), .Q(n3528) );
  INV15 U4720 ( .A(arg[29]), .Q(net713189) );
  NAND22 U4721 ( .A(n3973), .B(net715824), .Q(n3960) );
  CLKBU15 U4722 ( .A(n3574), .Q(n3578) );
  NAND22 U4723 ( .A(n3898), .B(net716390), .Q(n3956) );
  NOR42 U4724 ( .A(arg[31]), .B(arg[30]), .C(net719615), .D(net713189), .Q(
        n3579) );
  NAND24 U4725 ( .A(n4150), .B(n4149), .Q(n4214) );
  NAND21 U4726 ( .A(net723547), .B(net713055), .Q(net713152) );
  XNR22 U4727 ( .A(arg[23]), .B(n3063), .Q(n3632) );
  CLKBU15 U4728 ( .A(net715376), .Q(net715753) );
  NAND22 U4729 ( .A(n3747), .B(net712595), .Q(n3752) );
  BUF12 U4730 ( .A(N2561), .Q(n3542) );
  OAI212 U4731 ( .A(net718226), .B(n3263), .C(n4074), .Q(N2561) );
  INV12 U4732 ( .A(N2435), .Q(net715348) );
  OAI212 U4733 ( .A(net715739), .B(n4112), .C(n4111), .Q(n4276) );
  NAND24 U4734 ( .A(net713096), .B(net713167), .Q(net713146) );
  NAND24 U4735 ( .A(n4148), .B(n4147), .Q(n4212) );
  INV3 U4736 ( .A(N2688), .Q(n4134) );
  NAND28 U4737 ( .A(net720121), .B(net719603), .Q(net717814) );
  INV3 U4738 ( .A(N2689), .Q(n4132) );
  MUX24 U4739 ( .A(n3187), .B(N2861), .S(net720274), .Q(res_8_) );
  OAI212 U4740 ( .A(net721268), .B(n4116), .C(n4115), .Q(n4280) );
  NAND28 U4741 ( .A(n4014), .B(n4013), .Q(N2063) );
  NAND22 U4742 ( .A(net712605), .B(net723768), .Q(n3764) );
  INV6 U4743 ( .A(net712582), .Q(net712595) );
  AOI222 U4744 ( .A(n3981), .B(n3980), .C(n3979), .D(n3978), .Q(n3982) );
  INV6 U4745 ( .A(n3884), .Q(n3889) );
  INV6 U4746 ( .A(n4055), .Q(n4248) );
  OAI212 U4747 ( .A(net720894), .B(N2294), .C(n4070), .Q(n4071) );
  MUX21 U4748 ( .A(net715761), .B(N2955), .S(net711876), .Q(sqroot[5]) );
  MUX24 U4749 ( .A(n4219), .B(N2855), .S(net720274), .Q(res_2_) );
  INV12 U4750 ( .A(net716401), .Q(net716402) );
  INV0 U4751 ( .A(n3623), .Q(n3443) );
  NAND28 U4752 ( .A(n3450), .B(n3449), .Q(n3694) );
  NAND22 U4753 ( .A(arg[25]), .B(net718617), .Q(net718618) );
  NAND22 U4754 ( .A(net718604), .B(net718343), .Q(n3451) );
  NOR33 U4755 ( .A(n3460), .B(n3709), .C(net712716), .Q(n3712) );
  NAND22 U4756 ( .A(net712311), .B(n2913), .Q(n3462) );
  CLKIN6 U4757 ( .A(n3465), .Q(n3466) );
  NAND22 U4758 ( .A(net724837), .B(n2890), .Q(n3469) );
  NAND28 U4759 ( .A(n3469), .B(n3470), .Q(net712612) );
  XNR22 U4760 ( .A(net715614), .B(n3813), .Q(net712478) );
  INV6 U4761 ( .A(n3476), .Q(n3477) );
  NAND28 U4762 ( .A(n3479), .B(n3255), .Q(n3906) );
  NAND31 U4763 ( .A(net715700), .B(n3998), .C(n3997), .Q(n3999) );
  IMUX24 U4764 ( .A(n3795), .B(n3794), .S(net720787), .Q(n3796) );
  NAND34 U4765 ( .A(n3744), .B(n3745), .C(n3492), .Q(net712600) );
  INV6 U4766 ( .A(n3491), .Q(n3492) );
  INV1 U4767 ( .A(net712414), .Q(net718362) );
  NOR32 U4768 ( .A(net716172), .B(n3841), .C(n3840), .Q(n3842) );
  NAND22 U4769 ( .A(net712966), .B(net720967), .Q(n3496) );
  MUX22 U4770 ( .A(N1919), .B(N1790), .S(net715406), .Q(n3525) );
  NAND22 U4771 ( .A(N2499), .B(net718226), .Q(n3504) );
  NAND24 U4772 ( .A(n3503), .B(n3504), .Q(n3505) );
  NAND24 U4773 ( .A(n3615), .B(n3614), .Q(n3616) );
  XNR22 U4774 ( .A(n2947), .B(net712865), .Q(n3653) );
  AOI312 U4775 ( .A(n3946), .B(n3271), .C(n3945), .D(n2912), .Q(n3947) );
  OAI222 U4776 ( .A(N1784), .B(net715712), .C(n3923), .D(n3924), .Q(n3942) );
  NAND21 U4777 ( .A(N2876), .B(net719548), .Q(n4172) );
  NAND22 U4778 ( .A(N2854), .B(net715754), .Q(n4207) );
  NAND22 U4779 ( .A(N2874), .B(net722433), .Q(n4176) );
  NAND22 U4780 ( .A(N2877), .B(net719548), .Q(n4170) );
  INV3 U4781 ( .A(n3960), .Q(n3951) );
  NOR42 U4782 ( .A(n3731), .B(n3730), .C(n3250), .D(n3872), .Q(n3746) );
  OAI222 U4783 ( .A(N2291), .B(net718090), .C(n3441), .D(net715719), .Q(n4061)
         );
  OAI221 U4784 ( .A(n3885), .B(n3839), .C(n3863), .D(n3838), .Q(n3840) );
  OAI312 U4785 ( .A(n3678), .B(net712831), .C(n3669), .D(n3668), .Q(n3670) );
  XNR22 U4786 ( .A(arg[22]), .B(net715616), .Q(net712879) );
  XNR22 U4787 ( .A(n3244), .B(n3903), .Q(n4005) );
  OAI222 U4788 ( .A(net715719), .B(n3240), .C(N2285), .D(net718090), .Q(n4065)
         );
  XOR22 U4789 ( .A(n4004), .B(n4003), .Q(n3527) );
  NAND22 U4790 ( .A(N2284), .B(net718011), .Q(n3509) );
  NAND28 U4791 ( .A(n3508), .B(n3509), .Q(n3516) );
  AOI2111 U4792 ( .A(n4048), .B(net715767), .C(net715480), .D(net712145), .Q(
        n4036) );
  OAI212 U4793 ( .A(n3833), .B(n3543), .C(n3846), .Q(n3834) );
  CLKIN0 U4794 ( .A(net715710), .Q(net712990) );
  CLKIN2 U4795 ( .A(N2953), .Q(n3560) );
  CLKIN2 U4796 ( .A(N2952), .Q(n3559) );
  CLKIN2 U4797 ( .A(N2960), .Q(n3558) );
  CLKIN2 U4798 ( .A(N2962), .Q(n3561) );
  CLKIN2 U4799 ( .A(N2954), .Q(n3562) );
  CLKIN3 U4800 ( .A(arg[14]), .Q(net712454) );
  BUF2 U4801 ( .A(net715402), .Q(net715761) );
  MUX26 U4802 ( .A(n4254), .B(N2300), .S(net715717), .Q(n3521) );
  CLKIN0 U4803 ( .A(net715576), .Q(net715570) );
  AOI312 U4804 ( .A(n3567), .B(n3564), .C(n3966), .D(n3965), .Q(n3987) );
  INV3 U4805 ( .A(arg[15]), .Q(n3790) );
  MUX22 U4806 ( .A(n4262), .B(N2880), .S(net715754), .Q(res_27_) );
  MUX22 U4807 ( .A(n4261), .B(N2881), .S(net715753), .Q(res_28_) );
  INV3 U4808 ( .A(N1919), .Q(n4026) );
  BUF2 U4809 ( .A(n2927), .Q(net716101) );
  BUF2 U4810 ( .A(net715570), .Q(net715802) );
  BUF2 U4811 ( .A(net715478), .Q(net715782) );
  BUF2 U4812 ( .A(net715570), .Q(net715804) );
  BUF2 U4813 ( .A(net715478), .Q(net715783) );
  BUF2 U4814 ( .A(net715570), .Q(net715803) );
  BUF2 U4815 ( .A(net715478), .Q(net715781) );
  XOR22 U4816 ( .A(n3644), .B(n3643), .Q(n3724) );
  INV3 U4817 ( .A(net715610), .Q(net715606) );
  BUF2 U4818 ( .A(net675324), .Q(net715478) );
  BUF2 U4819 ( .A(net715769), .Q(net715776) );
  BUF2 U4820 ( .A(net715769), .Q(net715775) );
  AOI220 U4821 ( .A(n3817), .B(net712139), .C(n3819), .D(n3818), .Q(n3816) );
  AOI210 U4822 ( .A(net712899), .B(n3642), .C(net712901), .Q(n3644) );
  NAND20 U4823 ( .A(net712903), .B(net712904), .Q(n3642) );
  INV0 U4824 ( .A(net712902), .Q(net712901) );
  MUX21 U4825 ( .A(N2090), .B(n3534), .S(net715687), .Q(n4294) );
  MUX21 U4826 ( .A(net715816), .B(N2957), .S(net711876), .Q(sqroot[7]) );
  MUX21 U4827 ( .A(net720783), .B(N2958), .S(net711876), .Q(sqroot[8]) );
  MUX21 U4828 ( .A(net725733), .B(N2959), .S(net711876), .Q(sqroot[9]) );
  MUX21 U4829 ( .A(net715480), .B(N2964), .S(net711876), .Q(sqroot[14]) );
  MUX21 U4830 ( .A(net719772), .B(N2951), .S(net711876), .Q(sqroot[1]) );
  MUX21 U4831 ( .A(net721034), .B(N2950), .S(net711876), .Q(sqroot[0]) );
  IMUX21 U4832 ( .A(n4296), .B(N2280), .S(net715725), .Q(n4123) );
  MUX21 U4833 ( .A(N2088), .B(n3536), .S(net715687), .Q(n4296) );
  MUX21 U4834 ( .A(n4297), .B(N2279), .S(net723969), .Q(n3530) );
  MUX21 U4835 ( .A(N2086), .B(n3537), .S(net715687), .Q(n4298) );
  MUX21 U4836 ( .A(N1899), .B(arg[6]), .S(net715412), .Q(n3532) );
  MUX21 U4837 ( .A(N1900), .B(arg[7]), .S(net715412), .Q(n3533) );
  NAND22 U4838 ( .A(net713169), .B(net713170), .Q(n3594) );
  CLKIN3 U4839 ( .A(arg[29]), .Q(net713169) );
  MUX21 U4840 ( .A(N1898), .B(arg[5]), .S(net715412), .Q(n3534) );
  MUX21 U4841 ( .A(N1897), .B(arg[4]), .S(net715412), .Q(n3535) );
  MUX21 U4842 ( .A(N1896), .B(arg[3]), .S(net715412), .Q(n3536) );
  MUX21 U4843 ( .A(N1894), .B(arg[1]), .S(net715412), .Q(n3537) );
  MUX21 U4844 ( .A(N1895), .B(arg[2]), .S(net715412), .Q(n3538) );
  MUX21 U4845 ( .A(N1893), .B(arg[0]), .S(net715412), .Q(n3539) );
  LOGIC0 U4846 ( .Q(n4257) );
  LOGIC1 U4847 ( .Q(n4256) );
  NAND43 U4848 ( .A(n3957), .B(n3956), .C(n3955), .D(n3954), .Q(n3958) );
  NOR42 U4849 ( .A(n3917), .B(n3915), .C(n3506), .D(n3916), .Q(n3955) );
  XNR22 U4850 ( .A(net712993), .B(n3629), .Q(net712941) );
  NOR42 U4851 ( .A(n3267), .B(n3253), .C(net712634), .D(net712363), .Q(n3744)
         );
  NOR42 U4852 ( .A(net712816), .B(n3674), .C(n3661), .D(n3401), .Q(n3665) );
  AOI212 U4853 ( .A(net721041), .B(net726276), .C(n3557), .Q(n3556) );
  IMUX20 U4854 ( .A(net723435), .B(n3558), .S(net722521), .Q(sqroot[10]) );
  IMUX20 U4855 ( .A(net722422), .B(n3559), .S(net722521), .Q(sqroot[2]) );
  IMUX20 U4856 ( .A(net718067), .B(n3560), .S(net722521), .Q(sqroot[3]) );
  IMUX20 U4857 ( .A(net715576), .B(n3561), .S(net722521), .Q(sqroot[12]) );
  IMUX20 U4858 ( .A(n3578), .B(n3562), .S(net722521), .Q(sqroot[4]) );
  BUF2 U4859 ( .A(N1776), .Q(n3563) );
  XNR20 U4860 ( .A(net723637), .B(n3925), .Q(n3926) );
  BUF2 U4861 ( .A(n2884), .Q(net716222) );
  OAI211 U4862 ( .A(net712139), .B(n3230), .C(n4038), .Q(net712197) );
  CLKIN6 U4863 ( .A(n3870), .Q(N1786) );
  NOR32 U4864 ( .A(net712216), .B(net716172), .C(n3913), .Q(n3900) );
  NOR31 U4865 ( .A(n4004), .B(n2927), .C(n3990), .Q(n3991) );
  XNR22 U4866 ( .A(n3811), .B(net725181), .Q(n3950) );
  XNR22 U4867 ( .A(n3295), .B(n3693), .Q(n3812) );
  INV6 U4868 ( .A(n3986), .Q(n3572) );
  NAND34 U4869 ( .A(n3570), .B(n3571), .C(n3572), .Q(n3573) );
  NAND20 U4870 ( .A(n3960), .B(n3959), .Q(n3988) );
  XNR20 U4871 ( .A(n3543), .B(net715544), .Q(n3936) );
  XNR22 U4872 ( .A(n3313), .B(n3855), .Q(n3973) );
  XNR22 U4873 ( .A(n3257), .B(n3814), .Q(n3856) );
  NOR42 U4874 ( .A(n3461), .B(n3809), .C(n3810), .D(n3824), .Q(n3829) );
  NOR24 U4875 ( .A(n3793), .B(net712535), .Q(n3794) );
  XNR22 U4876 ( .A(net713043), .B(net713044), .Q(n3617) );
  INV6 U4877 ( .A(n3901), .Q(n3911) );
  OAI222 U4878 ( .A(N2287), .B(net718090), .C(n3324), .D(net719237), .Q(n4095)
         );
  MUX21 U4879 ( .A(N2085), .B(n3539), .S(n3578), .Q(n4299) );
  MUX21 U4880 ( .A(N2087), .B(n3538), .S(n3578), .Q(n4297) );
  MUX21 U4881 ( .A(N2089), .B(n3535), .S(n3578), .Q(n4295) );
  NAND28 U4882 ( .A(n4014), .B(n4013), .Q(net712208) );
  XNR22 U4883 ( .A(net723959), .B(net712433), .Q(N1780) );
  INV6 U4884 ( .A(n3588), .Q(n3590) );
  CLKIN3 U4885 ( .A(net715711), .Q(net675324) );
  CLKIN3 U4886 ( .A(n3592), .Q(n3581) );
  AOI2112 U4887 ( .A(n3581), .B(n3591), .C(n3580), .D(n3579), .Q(net713161) );
  AOI222 U4888 ( .A(n3280), .B(n3589), .C(n3582), .D(n3583), .Q(n3584) );
  OAI212 U4889 ( .A(n3585), .B(net713171), .C(n3584), .Q(net713181) );
  OAI212 U4890 ( .A(net715450), .B(net724021), .C(net715712), .Q(n3588) );
  OAI2112 U4891 ( .A(arg[26]), .B(n3017), .C(n3590), .D(arg[27]), .Q(net713149) );
  OAI212 U4892 ( .A(arg[29]), .B(arg[30]), .C(net713199), .Q(net713197) );
  CLKIN3 U4893 ( .A(net713186), .Q(net713196) );
  OAI222 U4894 ( .A(n3593), .B(net713189), .C(n3592), .D(n3591), .Q(net713167)
         );
  OAI2112 U4895 ( .A(n3595), .B(n3594), .C(net713166), .D(net715768), .Q(n3596) );
  CLKIN3 U4896 ( .A(arg[22]), .Q(net712963) );
  OAI212 U4897 ( .A(arg[26]), .B(net713157), .C(arg[27]), .Q(net713084) );
  NAND22 U4898 ( .A(net713099), .B(net721349), .Q(n3599) );
  OAI222 U4899 ( .A(arg[26]), .B(net713087), .C(net718490), .D(net713090), .Q(
        n3607) );
  NAND22 U4900 ( .A(n3604), .B(net713087), .Q(n3605) );
  XOR31 U4901 ( .A(n3610), .B(net715450), .C(n3609), .Q(n3611) );
  NAND22 U4902 ( .A(net712977), .B(net712976), .Q(net712970) );
  OAI212 U4903 ( .A(arg[25]), .B(net713055), .C(net715680), .Q(n3612) );
  OAI212 U4904 ( .A(net715680), .B(arg[25]), .C(net713051), .Q(n3614) );
  CLKIN3 U4905 ( .A(net713047), .Q(net713041) );
  NAND22 U4906 ( .A(net715480), .B(n3620), .Q(n3627) );
  NAND22 U4907 ( .A(n3627), .B(n3626), .Q(net713020) );
  NAND22 U4908 ( .A(n3623), .B(net715711), .Q(net713009) );
  NAND22 U4909 ( .A(net713020), .B(net713009), .Q(net713024) );
  CLKIN3 U4910 ( .A(arg[18]), .Q(net712793) );
  OAI212 U4911 ( .A(n3644), .B(n3643), .C(net712894), .Q(net712674) );
  OAI212 U4912 ( .A(net723702), .B(net712773), .C(net712774), .Q(net712766) );
  NAND22 U4913 ( .A(net712712), .B(net712760), .Q(n3689) );
  CLKIN3 U4914 ( .A(n3689), .Q(n3691) );
  XNR21 U4915 ( .A(n3691), .B(net712139), .Q(n3692) );
  NAND22 U4916 ( .A(net712454), .B(n3790), .Q(net712531) );
  OAI212 U4917 ( .A(net712754), .B(net712755), .C(net712730), .Q(n3697) );
  OAI212 U4918 ( .A(n3704), .B(n3713), .C(n3703), .Q(n3739) );
  CLKIN3 U4919 ( .A(n3732), .Q(n3733) );
  CLKIN3 U4920 ( .A(net712652), .Q(net712651) );
  OAI212 U4921 ( .A(net712642), .B(n3740), .C(net712644), .Q(n3743) );
  NAND22 U4922 ( .A(arg[16]), .B(net715544), .Q(net712505) );
  OAI212 U4923 ( .A(net712619), .B(net712620), .C(n3750), .Q(n3751) );
  OAI212 U4924 ( .A(net723577), .B(n3766), .C(n3268), .Q(n3767) );
  CLKIN3 U4925 ( .A(n3873), .Q(n3781) );
  NAND22 U4926 ( .A(n3781), .B(n3780), .Q(n3784) );
  OAI222 U4927 ( .A(arg[14]), .B(net712330), .C(arg[14]), .D(net712323), .Q(
        n3786) );
  OAI212 U4928 ( .A(net712139), .B(n3274), .C(n3832), .Q(n3809) );
  OAI212 U4929 ( .A(net712507), .B(n3484), .C(net719733), .Q(n3798) );
  CLKIN3 U4930 ( .A(n3799), .Q(n3807) );
  NAND22 U4931 ( .A(n3799), .B(net715608), .Q(n3802) );
  CLKIN3 U4932 ( .A(n3803), .Q(n3804) );
  AOI2112 U4933 ( .A(net723917), .B(n3807), .C(n3805), .D(n3806), .Q(n3808) );
  CLKIN3 U4934 ( .A(n3817), .Q(n3819) );
  AOI312 U4935 ( .A(n3822), .B(n3823), .C(n3821), .D(n3234), .Q(n3825) );
  OAI222 U4936 ( .A(n3826), .B(n3827), .C(n3824), .D(n3825), .Q(n3828) );
  NAND22 U4937 ( .A(net712323), .B(net712330), .Q(n3831) );
  CLKIN3 U4938 ( .A(n3831), .Q(n3925) );
  CLKIN3 U4939 ( .A(n3857), .Q(n3871) );
  CLKIN3 U4940 ( .A(n4000), .Q(n4004) );
  OAI212 U4941 ( .A(net712374), .B(n3881), .C(net712412), .Q(n3860) );
  OAI312 U4942 ( .A(n3865), .B(n3864), .C(n3863), .D(n3862), .Q(n3901) );
  XNR21 U4943 ( .A(n3207), .B(n3871), .Q(n4008) );
  CLKIN3 U4944 ( .A(n3874), .Q(n3876) );
  CLKIN3 U4945 ( .A(n3994), .Q(n3878) );
  NAND22 U4946 ( .A(n3996), .B(n3878), .Q(n3879) );
  OAI212 U4947 ( .A(n3882), .B(n2915), .C(n3881), .Q(n3884) );
  NAND22 U4948 ( .A(n3248), .B(n3889), .Q(n3892) );
  CLKIN3 U4949 ( .A(n3892), .Q(n3893) );
  OAI212 U4950 ( .A(net720567), .B(n3911), .C(net720570), .Q(n3913) );
  XNR21 U4951 ( .A(n3294), .B(n3907), .Q(n4002) );
  OAI312 U4952 ( .A(n4004), .B(n3909), .C(n3908), .D(n2889), .Q(N1793) );
  CLKIN3 U4953 ( .A(arg[8]), .Q(net712328) );
  CLKIN3 U4954 ( .A(arg[9]), .Q(n3918) );
  NAND22 U4955 ( .A(net712328), .B(n3918), .Q(n3919) );
  OAI222 U4956 ( .A(arg[10]), .B(arg[11]), .C(arg[11]), .D(n3919), .Q(n3921)
         );
  OAI212 U4957 ( .A(net720783), .B(n3935), .C(n3137), .Q(n3938) );
  CLKIN3 U4958 ( .A(arg[10]), .Q(n3961) );
  NAND22 U4959 ( .A(N1783), .B(net715678), .Q(n3980) );
  CLKIN3 U4960 ( .A(n3980), .Q(n3984) );
  OAI212 U4961 ( .A(n3984), .B(n3983), .C(n3982), .Q(n3985) );
  NAND22 U4962 ( .A(n3992), .B(n3996), .Q(n3993) );
  XNR21 U4963 ( .A(n3994), .B(n3993), .Q(n4226) );
  NAND22 U4964 ( .A(n4003), .B(n4000), .Q(n4001) );
  OAI222 U4965 ( .A(N1913), .B(net715416), .C(net725944), .D(net716390), .Q(
        n4048) );
  OAI212 U4966 ( .A(n4018), .B(n4017), .C(n4021), .Q(n4019) );
  AOI212 U4967 ( .A(net712171), .B(n4023), .C(n4022), .Q(net712169) );
  OAI222 U4968 ( .A(net715759), .B(n3192), .C(n4029), .D(n4028), .Q(net712151)
         );
  OAI222 U4969 ( .A(n4030), .B(n4031), .C(net715769), .D(n4048), .Q(n4032) );
  AOI212 U4970 ( .A(n4037), .B(N1974), .C(n4036), .Q(net712126) );
  OAI222 U4971 ( .A(n4041), .B(n4040), .C(n3341), .D(net715788), .Q(n4042) );
  CLKIN3 U4972 ( .A(n4043), .Q(N1987) );
  CLKIN3 U4973 ( .A(n4044), .Q(N1986) );
  CLKIN3 U4974 ( .A(n4045), .Q(N1983) );
  CLKIN3 U4975 ( .A(n4046), .Q(N1981) );
  CLKIN3 U4976 ( .A(n4047), .Q(N1980) );
  NAND22 U4977 ( .A(N2114), .B(n3576), .Q(n4049) );
  OAI222 U4978 ( .A(n3237), .B(n4056), .C(net715717), .D(n3237), .Q(n4230) );
  OAI222 U4979 ( .A(net722482), .B(n4059), .C(n4058), .D(n4059), .Q(n4227) );
  OAI222 U4980 ( .A(n4060), .B(n3306), .C(n3306), .D(net722482), .Q(n4228) );
  OAI222 U4981 ( .A(N2290), .B(net718067), .C(net715719), .D(n3522), .Q(n4090)
         );
  OAI222 U4982 ( .A(net715719), .B(n3238), .C(N2286), .D(net718090), .Q(n4097)
         );
  OAI222 U4983 ( .A(N2283), .B(net719234), .C(net715719), .D(n4293), .Q(n4099)
         );
  OAI222 U4984 ( .A(net715719), .B(n4294), .C(N2282), .D(net718090), .Q(n4066)
         );
  CLKIN3 U4985 ( .A(n4123), .Q(n4235) );
  CLKIN3 U4986 ( .A(n4125), .Q(n4234) );
  OAI212 U4987 ( .A(N2295), .B(net718067), .C(n4068), .Q(n4069) );
  OAI212 U4988 ( .A(net719234), .B(N2293), .C(n3417), .Q(n4089) );
  OAI212 U4989 ( .A(net719306), .B(n4079), .C(n4078), .Q(N2557) );
  OAI212 U4990 ( .A(net719306), .B(n4084), .C(n4083), .Q(N2553) );
  OAI212 U4991 ( .A(net717907), .B(n4093), .C(n4092), .Q(N2543) );
  OAI212 U4992 ( .A(net718129), .B(n3357), .C(n4094), .Q(N2542) );
  OAI212 U4993 ( .A(net723620), .B(n3301), .C(n4096), .Q(N2541) );
  NAND22 U4994 ( .A(N2691), .B(net722561), .Q(n4127) );
  NAND22 U4995 ( .A(n3505), .B(net715360), .Q(n4128) );
  NAND22 U4996 ( .A(n4127), .B(n4128), .Q(n4259) );
  NAND22 U4997 ( .A(N2690), .B(net722561), .Q(n4129) );
  NAND22 U4998 ( .A(n3542), .B(net719771), .Q(n4130) );
  NAND22 U4999 ( .A(n4129), .B(n4130), .Q(n4260) );
  NAND22 U5000 ( .A(N2560), .B(net715360), .Q(n4131) );
  NAND22 U5001 ( .A(n3454), .B(net722560), .Q(n4136) );
  NAND22 U5002 ( .A(n4137), .B(n4138), .Q(n4264) );
  NAND22 U5003 ( .A(n3517), .B(net719771), .Q(n4141) );
  NAND22 U5004 ( .A(N2681), .B(net722561), .Q(n4148) );
  OAI212 U5005 ( .A(net722561), .B(n3395), .C(n4105), .Q(n4272) );
  OAI212 U5006 ( .A(net721268), .B(n4108), .C(n4107), .Q(n4273) );
  OAI212 U5007 ( .A(net715739), .B(n4114), .C(n4113), .Q(n4277) );
  OAI222 U5008 ( .A(net719447), .B(n4154), .C(net715739), .D(n4153), .Q(n4223)
         );
  OAI212 U5009 ( .A(net721268), .B(n4118), .C(n4117), .Q(n4281) );
  OAI212 U5010 ( .A(net721268), .B(n3266), .C(n4121), .Q(n4283) );
  NAND22 U5011 ( .A(net717664), .B(N2665), .Q(net711939) );
  OAI212 U5012 ( .A(net721268), .B(n4123), .C(n4122), .Q(n4284) );
  NAND22 U5013 ( .A(net717664), .B(N2663), .Q(n4157) );
  NAND22 U5014 ( .A(n4157), .B(n4158), .Q(n4219) );
  NAND22 U5015 ( .A(net718162), .B(N2662), .Q(n4124) );
  OAI212 U5016 ( .A(net715739), .B(n4125), .C(n4124), .Q(n4286) );
  CLKIN3 U5017 ( .A(N2661), .Q(n4126) );
  CLKIN3 U5018 ( .A(n4209), .Q(n4287) );
  NAND22 U5019 ( .A(n4128), .B(n4127), .Q(n4216) );
  NAND22 U5020 ( .A(n4130), .B(n4129), .Q(n4224) );
  OAI212 U5021 ( .A(net715360), .B(n4132), .C(n4131), .Q(n4261) );
  OAI212 U5022 ( .A(net715360), .B(n4134), .C(n4133), .Q(n4262) );
  NAND22 U5023 ( .A(n4136), .B(n4135), .Q(n4218) );
  NAND22 U5024 ( .A(n4140), .B(n4139), .Q(n4213) );
  NAND22 U5025 ( .A(n4142), .B(n4141), .Q(n4215) );
  OAI212 U5026 ( .A(net715360), .B(n4152), .C(n4151), .Q(n4222) );
  OAI222 U5027 ( .A(net719447), .B(n4154), .C(net715739), .D(n4153), .Q(n4278)
         );
  CLKIN3 U5028 ( .A(n4216), .Q(n4163) );
  OAI212 U5029 ( .A(net721034), .B(n4163), .C(n4162), .Q(res_30_) );
  CLKIN3 U5030 ( .A(n4224), .Q(n4165) );
  OAI212 U5031 ( .A(net719548), .B(n4165), .C(n4164), .Q(res_29_) );
  CLKIN3 U5032 ( .A(n4218), .Q(n4167) );
  OAI212 U5033 ( .A(net719548), .B(n4167), .C(n4166), .Q(res_26_) );
  CLKIN3 U5034 ( .A(n4221), .Q(n4169) );
  CLKIN3 U5035 ( .A(n4213), .Q(n4171) );
  OAI212 U5036 ( .A(net719548), .B(n4171), .C(n4170), .Q(res_24_) );
  NAND22 U5037 ( .A(N2875), .B(net721034), .Q(n4174) );
  OAI212 U5038 ( .A(net721034), .B(n4177), .C(n4176), .Q(res_21_) );
  CLKIN3 U5039 ( .A(n4212), .Q(n4179) );
  OAI212 U5040 ( .A(net719548), .B(n4179), .C(n4178), .Q(res_20_) );
  CLKIN3 U5041 ( .A(n4214), .Q(n4181) );
  NAND22 U5042 ( .A(N2872), .B(net719548), .Q(n4180) );
  OAI212 U5043 ( .A(net715754), .B(n4186), .C(n4185), .Q(res_17_) );
  OAI212 U5044 ( .A(net715754), .B(n4188), .C(n4187), .Q(res_15_) );
  NAND22 U5045 ( .A(N2867), .B(net715754), .Q(n4189) );
  OAI212 U5046 ( .A(net722433), .B(n4190), .C(n4189), .Q(res_14_) );
  OAI212 U5047 ( .A(net711901), .B(net715753), .C(n4191), .Q(res_13_) );
  OAI212 U5048 ( .A(net715753), .B(n4193), .C(n4192), .Q(res_12_) );
  CLKIN3 U5049 ( .A(n3544), .Q(n4201) );
  OAI212 U5050 ( .A(n4203), .B(net720325), .C(n4202), .Q(res_6_) );
  OAI212 U5051 ( .A(net715753), .B(n4205), .C(n4204), .Q(res_5_) );
  OAI212 U5052 ( .A(net715754), .B(n4208), .C(n4207), .Q(res_1_) );
  XNR21 U5053 ( .A(n4209), .B(net715753), .Q(res_0_) );
endmodule

