
module sqroot_seq_NBITS32_DW01_inc_1 ( A, SUM );
  input [31:0] A;
  output [31:0] SUM;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n17,
         n18, n19, n20, n22, n23, n24, n25, n26, n28, n29, n30, n31, n33, n34,
         n35, n36, n37, n40, n41, n42, n45, n46, n47, n49, n50, n52, n53, n54,
         n55, n57, n58, n59, n60, n61, n64, n65, n66, n69, n70, n71, n72, n74,
         n76, n77, n78, n81, n82, n83, n84, n88, n89, n91, n93, n94, n95, n97,
         n98, n99, n100, n102, n103, n104, n105, n106, n109, n110, n111, n114,
         n115, n116, n117, n119, n121, n122, n123, n126, n127, n128, n129,
         n134, n137, n138, n139, n140, n142, n143, n144, n146, n147, n148,
         n149, n152, n153, n156, n157, n158, n159, n161, n162, n165, n166,
         n238, n239, n240, n241;

  NAND20 U204 ( .A(n149), .B(A[6]), .Q(n144) );
  NOR21 U205 ( .A(n50), .B(n60), .Q(n49) );
  NAND22 U206 ( .A(A[20]), .B(A[21]), .Q(n60) );
  NAND24 U207 ( .A(A[16]), .B(A[17]), .Q(n84) );
  INV8 U208 ( .A(n238), .Q(n239) );
  INV3 U209 ( .A(n71), .Q(n72) );
  XOR21 U210 ( .A(n88), .B(n89), .Q(SUM[17]) );
  XNR21 U211 ( .A(n91), .B(n239), .Q(SUM[16]) );
  NOR23 U212 ( .A(n95), .B(n105), .Q(n94) );
  NOR22 U213 ( .A(n140), .B(n148), .Q(n139) );
  NAND23 U214 ( .A(A[8]), .B(A[9]), .Q(n129) );
  NAND22 U215 ( .A(n241), .B(n83), .Q(n82) );
  INV3 U216 ( .A(n116), .Q(n117) );
  NOR23 U217 ( .A(n138), .B(n93), .Q(n2) );
  XOR21 U218 ( .A(n102), .B(n103), .Q(SUM[14]) );
  INV3 U219 ( .A(n166), .Q(n165) );
  NAND23 U220 ( .A(A[1]), .B(A[0]), .Q(n166) );
  NOR23 U221 ( .A(n26), .B(n36), .Q(n4) );
  NAND22 U222 ( .A(A[26]), .B(A[27]), .Q(n26) );
  NOR20 U223 ( .A(n60), .B(n72), .Q(n59) );
  INV6 U224 ( .A(n138), .Q(n137) );
  NAND22 U225 ( .A(n239), .B(n78), .Q(n77) );
  INV3 U226 ( .A(n148), .Q(n149) );
  NOR21 U227 ( .A(n144), .B(n157), .Q(n143) );
  INV1 U228 ( .A(A[12]), .Q(n114) );
  NAND22 U229 ( .A(A[4]), .B(A[5]), .Q(n148) );
  XOR21 U230 ( .A(A[8]), .B(n137), .Q(SUM[8]) );
  XOR21 U231 ( .A(n76), .B(n77), .Q(SUM[19]) );
  CLKIN6 U232 ( .A(n158), .Q(n157) );
  XNR21 U233 ( .A(n152), .B(n153), .Q(SUM[5]) );
  NAND22 U234 ( .A(A[6]), .B(A[7]), .Q(n140) );
  NAND21 U235 ( .A(n42), .B(n241), .Q(n41) );
  NOR20 U236 ( .A(n45), .B(n3), .Q(n42) );
  INV6 U237 ( .A(n240), .Q(n241) );
  NAND28 U238 ( .A(n139), .B(n158), .Q(n138) );
  XOR20 U239 ( .A(n161), .B(n162), .Q(SUM[3]) );
  NAND20 U240 ( .A(n165), .B(A[2]), .Q(n162) );
  XOR21 U241 ( .A(n81), .B(n82), .Q(SUM[18]) );
  NAND22 U242 ( .A(n241), .B(n47), .Q(n46) );
  XOR21 U243 ( .A(n69), .B(n70), .Q(SUM[20]) );
  NAND23 U244 ( .A(A[10]), .B(A[11]), .Q(n119) );
  NOR24 U245 ( .A(n119), .B(n129), .Q(n116) );
  NAND22 U246 ( .A(n116), .B(n94), .Q(n93) );
  NAND22 U247 ( .A(n137), .B(n116), .Q(n115) );
  NOR24 U248 ( .A(n166), .B(n159), .Q(n158) );
  NAND22 U249 ( .A(n239), .B(A[16]), .Q(n89) );
  NAND22 U250 ( .A(n30), .B(n241), .Q(n29) );
  NAND22 U251 ( .A(n137), .B(n123), .Q(n122) );
  NAND22 U252 ( .A(A[2]), .B(A[3]), .Q(n159) );
  NAND22 U253 ( .A(n137), .B(n128), .Q(n127) );
  CLKIN6 U254 ( .A(n2), .Q(n238) );
  XOR21 U255 ( .A(n114), .B(n115), .Q(SUM[12]) );
  NAND21 U256 ( .A(n24), .B(n239), .Q(n23) );
  NAND22 U257 ( .A(n239), .B(n66), .Q(n65) );
  NAND21 U258 ( .A(n35), .B(n239), .Q(n34) );
  NAND22 U259 ( .A(n99), .B(n137), .Q(n98) );
  NOR20 U260 ( .A(n100), .B(n117), .Q(n99) );
  NAND22 U261 ( .A(n241), .B(n71), .Q(n70) );
  XOR21 U262 ( .A(n121), .B(n122), .Q(SUM[11]) );
  NAND21 U263 ( .A(n111), .B(n137), .Q(n110) );
  NOR20 U264 ( .A(n114), .B(n117), .Q(n111) );
  NAND22 U265 ( .A(n137), .B(A[8]), .Q(n134) );
  XOR21 U266 ( .A(n64), .B(n65), .Q(SUM[21]) );
  NAND21 U267 ( .A(n104), .B(n137), .Q(n103) );
  NAND22 U268 ( .A(n239), .B(n54), .Q(n53) );
  NOR21 U269 ( .A(n55), .B(n72), .Q(n54) );
  NAND21 U270 ( .A(A[18]), .B(A[19]), .Q(n74) );
  NAND22 U271 ( .A(n241), .B(n59), .Q(n58) );
  INV0 U272 ( .A(n36), .Q(n37) );
  NAND22 U273 ( .A(A[12]), .B(A[13]), .Q(n105) );
  NAND21 U274 ( .A(A[24]), .B(A[25]), .Q(n36) );
  NAND22 U275 ( .A(n37), .B(A[26]), .Q(n31) );
  NOR21 U276 ( .A(n126), .B(n129), .Q(n123) );
  XOR21 U277 ( .A(n22), .B(n23), .Q(SUM[28]) );
  XOR21 U278 ( .A(n29), .B(n28), .Q(SUM[27]) );
  XOR21 U279 ( .A(n109), .B(n110), .Q(SUM[13]) );
  XOR21 U280 ( .A(n33), .B(n34), .Q(SUM[26]) );
  XOR20 U281 ( .A(n126), .B(n127), .Q(SUM[10]) );
  XOR21 U282 ( .A(n40), .B(n41), .Q(SUM[25]) );
  XOR21 U283 ( .A(n52), .B(n53), .Q(SUM[23]) );
  NAND22 U284 ( .A(A[14]), .B(A[15]), .Q(n95) );
  NAND20 U285 ( .A(A[28]), .B(A[29]), .Q(n15) );
  CLKIN6 U286 ( .A(n2), .Q(n240) );
  CLKIN0 U287 ( .A(A[15]), .Q(n97) );
  NOR20 U288 ( .A(n148), .B(n157), .Q(n147) );
  XOR20 U289 ( .A(n156), .B(n157), .Q(SUM[4]) );
  NOR20 U290 ( .A(n105), .B(n117), .Q(n104) );
  XNR21 U291 ( .A(A[9]), .B(n134), .Q(SUM[9]) );
  XOR20 U292 ( .A(n57), .B(n58), .Q(SUM[22]) );
  NAND24 U293 ( .A(n71), .B(n49), .Q(n3) );
  NAND22 U294 ( .A(A[22]), .B(A[23]), .Q(n50) );
  INV0 U295 ( .A(A[0]), .Q(SUM[0]) );
  XNR21 U296 ( .A(n146), .B(n147), .Q(SUM[6]) );
  XOR20 U297 ( .A(n45), .B(n46), .Q(SUM[24]) );
  CLKIN0 U298 ( .A(A[18]), .Q(n81) );
  CLKIN0 U299 ( .A(A[16]), .Q(n91) );
  CLKIN0 U300 ( .A(A[20]), .Q(n69) );
  NOR20 U301 ( .A(n20), .B(n3), .Q(n19) );
  NAND20 U302 ( .A(n4), .B(A[28]), .Q(n20) );
  CLKIN0 U303 ( .A(A[17]), .Q(n88) );
  CLKIN0 U304 ( .A(A[13]), .Q(n109) );
  CLKIN0 U305 ( .A(A[14]), .Q(n102) );
  CLKIN0 U306 ( .A(A[26]), .Q(n33) );
  XOR20 U307 ( .A(n17), .B(n18), .Q(SUM[29]) );
  XOR21 U308 ( .A(n10), .B(n11), .Q(SUM[30]) );
  INV0 U309 ( .A(n105), .Q(n106) );
  INV0 U310 ( .A(n60), .Q(n61) );
  CLKIN0 U311 ( .A(A[27]), .Q(n28) );
  INV0 U312 ( .A(A[29]), .Q(n17) );
  NOR21 U313 ( .A(n156), .B(n157), .Q(n153) );
  CLKIN0 U314 ( .A(A[10]), .Q(n126) );
  NOR21 U315 ( .A(n25), .B(n3), .Q(n24) );
  INV3 U316 ( .A(n4), .Q(n25) );
  NOR21 U317 ( .A(n36), .B(n3), .Q(n35) );
  NAND20 U318 ( .A(n12), .B(n239), .Q(n11) );
  NOR21 U319 ( .A(n13), .B(n3), .Q(n12) );
  NAND22 U320 ( .A(n4), .B(n14), .Q(n13) );
  INV3 U321 ( .A(n15), .Q(n14) );
  NOR21 U322 ( .A(n81), .B(n84), .Q(n78) );
  INV3 U323 ( .A(n129), .Q(n128) );
  NOR20 U324 ( .A(n69), .B(n72), .Q(n66) );
  INV3 U325 ( .A(n3), .Q(n47) );
  INV3 U326 ( .A(n84), .Q(n83) );
  NAND20 U327 ( .A(n7), .B(n241), .Q(n6) );
  NOR21 U328 ( .A(n8), .B(n3), .Q(n7) );
  NAND22 U329 ( .A(n4), .B(n9), .Q(n8) );
  NOR21 U330 ( .A(n10), .B(n15), .Q(n9) );
  XOR21 U331 ( .A(n5), .B(n6), .Q(SUM[31]) );
  XOR21 U332 ( .A(n97), .B(n98), .Q(SUM[15]) );
  NOR22 U333 ( .A(n74), .B(n84), .Q(n71) );
  XNR21 U334 ( .A(n142), .B(n143), .Q(SUM[7]) );
  CLKIN0 U335 ( .A(A[24]), .Q(n45) );
  INV0 U336 ( .A(A[28]), .Q(n22) );
  INV0 U337 ( .A(A[21]), .Q(n64) );
  INV0 U338 ( .A(A[25]), .Q(n40) );
  INV0 U339 ( .A(A[22]), .Q(n57) );
  INV0 U340 ( .A(A[19]), .Q(n76) );
  INV0 U341 ( .A(A[23]), .Q(n52) );
  XOR20 U342 ( .A(A[2]), .B(n165), .Q(SUM[2]) );
  XOR20 U343 ( .A(A[0]), .B(A[1]), .Q(SUM[1]) );
  NOR21 U344 ( .A(n31), .B(n3), .Q(n30) );
  NAND20 U345 ( .A(n19), .B(n241), .Q(n18) );
  NAND20 U346 ( .A(n106), .B(A[14]), .Q(n100) );
  NAND20 U347 ( .A(n61), .B(A[22]), .Q(n55) );
  INV3 U348 ( .A(A[30]), .Q(n10) );
  INV3 U349 ( .A(A[31]), .Q(n5) );
  INV1 U350 ( .A(A[4]), .Q(n156) );
  INV0 U351 ( .A(A[7]), .Q(n142) );
  INV0 U352 ( .A(A[11]), .Q(n121) );
  INV0 U353 ( .A(A[5]), .Q(n152) );
  INV0 U354 ( .A(A[3]), .Q(n161) );
  INV0 U355 ( .A(A[6]), .Q(n146) );
endmodule


module sqroot_seq_NBITS32_DW_cmp_5 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181;

  OAI212 U1 ( .A(n1), .B(n21), .C(n2), .Q(GE_LT_GT_LE) );
  OAI212 U24 ( .A(n39), .B(n24), .C(n25), .Q(n23) );
  AOI212 U26 ( .A(n33), .B(n26), .C(n27), .Q(n25) );
  OAI212 U28 ( .A(n31), .B(n28), .C(n29), .Q(n27) );
  AOI212 U40 ( .A(n47), .B(n40), .C(n41), .Q(n39) );
  OAI212 U42 ( .A(n45), .B(n42), .C(n43), .Q(n41) );
  OAI212 U48 ( .A(n51), .B(n48), .C(n49), .Q(n47) );
  OAI212 U53 ( .A(n75), .B(n53), .C(n54), .Q(n52) );
  OAI212 U57 ( .A(n60), .B(n57), .C(n58), .Q(n56) );
  OAI212 U63 ( .A(n63), .B(n66), .C(n64), .Q(n62) );
  AOI212 U76 ( .A(n98), .B(n76), .C(n77), .Q(n75) );
  OAI212 U78 ( .A(n89), .B(n78), .C(n79), .Q(n77) );
  OAI212 U99 ( .A(n99), .B(n109), .C(n100), .Q(n98) );
  OAI212 U112 ( .A(n115), .B(n112), .C(n113), .Q(n111) );
  OAI212 U117 ( .A(n117), .B(n127), .C(n118), .Q(n116) );
  OAI212 U133 ( .A(n143), .B(n133), .C(n134), .Q(n132) );
  AOI212 U187 ( .A(n132), .B(n128), .C(n129), .Q(n127) );
  NAND23 U188 ( .A(n26), .B(n32), .Q(n24) );
  NOR22 U189 ( .A(n180), .B(B[30]), .Q(n9) );
  NOR23 U190 ( .A(n174), .B(B[24]), .Q(n36) );
  NAND22 U191 ( .A(B[12]), .B(n162), .Q(n93) );
  INV3 U192 ( .A(n82), .Q(n80) );
  NOR22 U193 ( .A(n42), .B(n44), .Q(n40) );
  AOI211 U194 ( .A(n62), .B(n55), .C(n56), .Q(n54) );
  CLKIN3 U195 ( .A(A[16]), .Q(n166) );
  NOR24 U196 ( .A(n177), .B(B[27]), .Q(n28) );
  NOR23 U197 ( .A(n164), .B(B[14]), .Q(n82) );
  NAND23 U198 ( .A(n84), .B(n80), .Q(n78) );
  NAND22 U199 ( .A(B[11]), .B(n161), .Q(n97) );
  NAND22 U200 ( .A(B[14]), .B(n164), .Q(n83) );
  NOR21 U201 ( .A(n171), .B(B[21]), .Q(n48) );
  NAND21 U202 ( .A(B[24]), .B(n174), .Q(n37) );
  NOR22 U203 ( .A(n88), .B(n78), .Q(n76) );
  NOR21 U204 ( .A(n161), .B(B[11]), .Q(n96) );
  NAND21 U205 ( .A(B[18]), .B(n168), .Q(n60) );
  NOR21 U206 ( .A(n65), .B(n63), .Q(n61) );
  NOR21 U207 ( .A(n57), .B(n59), .Q(n55) );
  NOR22 U208 ( .A(n168), .B(B[18]), .Q(n59) );
  NOR21 U209 ( .A(n9), .B(n11), .Q(n7) );
  NAND22 U210 ( .A(n55), .B(n61), .Q(n53) );
  NOR22 U211 ( .A(n165), .B(B[15]), .Q(n73) );
  CLKIN3 U212 ( .A(n125), .Q(n123) );
  NAND22 U213 ( .A(B[15]), .B(n165), .Q(n74) );
  INV2 U214 ( .A(n74), .Q(n72) );
  NOR23 U215 ( .A(n173), .B(B[23]), .Q(n42) );
  NAND20 U216 ( .A(B[23]), .B(n173), .Q(n43) );
  NOR22 U217 ( .A(n175), .B(B[25]), .Q(n34) );
  NOR22 U218 ( .A(n36), .B(n34), .Q(n32) );
  NAND22 U219 ( .A(B[22]), .B(n172), .Q(n45) );
  OAI212 U220 ( .A(n9), .B(n12), .C(n10), .Q(n8) );
  AOI212 U221 ( .A(n13), .B(n18), .C(n14), .Q(n12) );
  INV2 U222 ( .A(n73), .Q(n71) );
  NAND22 U223 ( .A(B[17]), .B(n167), .Q(n64) );
  NOR22 U224 ( .A(n167), .B(B[17]), .Q(n63) );
  NAND20 U225 ( .A(B[19]), .B(n169), .Q(n58) );
  NOR22 U226 ( .A(n38), .B(n24), .Q(n22) );
  NOR22 U227 ( .A(n155), .B(B[5]), .Q(n125) );
  CLKIN0 U228 ( .A(A[20]), .Q(n170) );
  AOI212 U229 ( .A(n90), .B(n95), .C(n91), .Q(n89) );
  INV6 U230 ( .A(n92), .Q(n90) );
  INV0 U231 ( .A(A[13]), .Q(n163) );
  CLKIN0 U232 ( .A(A[6]), .Q(n156) );
  AOI212 U233 ( .A(n80), .B(n85), .C(n81), .Q(n79) );
  OAI211 U234 ( .A(n37), .B(n34), .C(n35), .Q(n33) );
  NAND20 U235 ( .A(B[25]), .B(n175), .Q(n35) );
  CLKIN3 U236 ( .A(A[12]), .Q(n162) );
  AOI212 U237 ( .A(n110), .B(n116), .C(n111), .Q(n109) );
  NOR24 U238 ( .A(n166), .B(B[16]), .Q(n69) );
  CLKIN6 U239 ( .A(n69), .Q(n67) );
  NOR22 U240 ( .A(n172), .B(B[22]), .Q(n44) );
  NOR21 U241 ( .A(n170), .B(B[20]), .Q(n50) );
  NOR24 U242 ( .A(n162), .B(B[12]), .Q(n92) );
  NOR23 U243 ( .A(n28), .B(n30), .Q(n26) );
  NOR22 U244 ( .A(n176), .B(B[26]), .Q(n30) );
  NAND22 U245 ( .A(n67), .B(n71), .Q(n65) );
  NOR22 U246 ( .A(n169), .B(B[19]), .Q(n57) );
  NAND22 U247 ( .A(B[27]), .B(n177), .Q(n29) );
  NAND22 U248 ( .A(n17), .B(n13), .Q(n11) );
  INV0 U249 ( .A(A[31]), .Q(n181) );
  NAND21 U250 ( .A(B[26]), .B(n176), .Q(n31) );
  AOI212 U251 ( .A(n22), .B(n52), .C(n23), .Q(n21) );
  AOI212 U252 ( .A(n8), .B(n3), .C(n4), .Q(n2) );
  INV2 U253 ( .A(n6), .Q(n4) );
  INV2 U254 ( .A(n104), .Q(n102) );
  CLKIN3 U255 ( .A(n121), .Q(n119) );
  AOI212 U256 ( .A(n67), .B(n72), .C(n68), .Q(n66) );
  NAND22 U257 ( .A(n94), .B(n90), .Q(n88) );
  INV2 U258 ( .A(n96), .Q(n94) );
  NAND20 U259 ( .A(B[21]), .B(n171), .Q(n49) );
  NAND21 U260 ( .A(B[4]), .B(n154), .Q(n131) );
  INV2 U261 ( .A(n19), .Q(n17) );
  NOR20 U262 ( .A(n178), .B(B[28]), .Q(n19) );
  NAND20 U263 ( .A(B[29]), .B(n179), .Q(n16) );
  INV0 U264 ( .A(A[2]), .Q(n152) );
  INV0 U265 ( .A(A[1]), .Q(n151) );
  INV0 U266 ( .A(A[29]), .Q(n179) );
  INV0 U267 ( .A(A[7]), .Q(n157) );
  INV2 U268 ( .A(n103), .Q(n101) );
  NOR21 U269 ( .A(n160), .B(B[10]), .Q(n103) );
  INV2 U270 ( .A(n107), .Q(n105) );
  INV2 U271 ( .A(n108), .Q(n106) );
  INV0 U272 ( .A(A[9]), .Q(n159) );
  CLKIN3 U273 ( .A(n130), .Q(n128) );
  CLKIN3 U274 ( .A(n141), .Q(n139) );
  NAND21 U275 ( .A(B[28]), .B(n178), .Q(n20) );
  INV2 U276 ( .A(n93), .Q(n91) );
  NAND21 U277 ( .A(B[3]), .B(n153), .Q(n138) );
  CLKIN2 U278 ( .A(n146), .Q(n144) );
  CLKIN3 U279 ( .A(n142), .Q(n140) );
  NAND21 U280 ( .A(B[2]), .B(n152), .Q(n142) );
  NAND21 U281 ( .A(B[6]), .B(n156), .Q(n122) );
  NAND22 U282 ( .A(n7), .B(n3), .Q(n1) );
  AOI211 U283 ( .A(n119), .B(n124), .C(n120), .Q(n118) );
  NAND22 U284 ( .A(n119), .B(n123), .Q(n117) );
  INV3 U285 ( .A(n83), .Q(n81) );
  AOI211 U286 ( .A(n101), .B(n106), .C(n102), .Q(n100) );
  NAND22 U287 ( .A(n101), .B(n105), .Q(n99) );
  AOI211 U288 ( .A(n144), .B(n148), .C(n145), .Q(n143) );
  NAND22 U289 ( .A(n135), .B(n139), .Q(n133) );
  AOI211 U290 ( .A(n135), .B(n140), .C(n136), .Q(n134) );
  INV3 U291 ( .A(n5), .Q(n3) );
  NOR21 U292 ( .A(n181), .B(B[31]), .Q(n5) );
  NAND21 U293 ( .A(B[31]), .B(n181), .Q(n6) );
  NOR22 U294 ( .A(n158), .B(B[8]), .Q(n112) );
  NAND22 U295 ( .A(B[7]), .B(n157), .Q(n115) );
  NAND20 U296 ( .A(B[8]), .B(n158), .Q(n113) );
  NOR21 U297 ( .A(n156), .B(B[6]), .Q(n121) );
  NAND21 U298 ( .A(B[20]), .B(n170), .Q(n51) );
  INV3 U299 ( .A(n16), .Q(n14) );
  INV3 U300 ( .A(n137), .Q(n135) );
  NOR21 U301 ( .A(n153), .B(B[3]), .Q(n137) );
  NOR21 U302 ( .A(n152), .B(B[2]), .Q(n141) );
  INV3 U303 ( .A(n122), .Q(n120) );
  NOR21 U304 ( .A(n114), .B(n112), .Q(n110) );
  NOR21 U305 ( .A(n157), .B(B[7]), .Q(n114) );
  INV3 U306 ( .A(n15), .Q(n13) );
  NOR21 U307 ( .A(n179), .B(B[29]), .Q(n15) );
  INV3 U308 ( .A(n86), .Q(n84) );
  NOR21 U309 ( .A(n163), .B(B[13]), .Q(n86) );
  NOR20 U310 ( .A(n159), .B(B[9]), .Q(n107) );
  INV3 U311 ( .A(n126), .Q(n124) );
  NAND22 U312 ( .A(B[5]), .B(n155), .Q(n126) );
  NAND22 U313 ( .A(n46), .B(n40), .Q(n38) );
  NOR21 U314 ( .A(n48), .B(n50), .Q(n46) );
  NOR21 U315 ( .A(n154), .B(B[4]), .Q(n130) );
  NAND20 U316 ( .A(B[9]), .B(n159), .Q(n108) );
  INV3 U317 ( .A(n131), .Q(n129) );
  NAND20 U318 ( .A(B[10]), .B(n160), .Q(n104) );
  INV3 U319 ( .A(n138), .Q(n136) );
  INV3 U320 ( .A(n147), .Q(n145) );
  NAND22 U321 ( .A(B[1]), .B(n151), .Q(n147) );
  INV3 U322 ( .A(n87), .Q(n85) );
  NOR21 U323 ( .A(n151), .B(B[1]), .Q(n146) );
  INV3 U324 ( .A(n97), .Q(n95) );
  INV3 U325 ( .A(n20), .Q(n18) );
  INV3 U326 ( .A(n70), .Q(n68) );
  NAND22 U327 ( .A(B[16]), .B(n166), .Q(n70) );
  INV3 U328 ( .A(A[10]), .Q(n160) );
  INV0 U329 ( .A(A[4]), .Q(n154) );
  INV0 U330 ( .A(A[28]), .Q(n178) );
  INV3 U331 ( .A(A[25]), .Q(n175) );
  CLKIN0 U332 ( .A(A[3]), .Q(n153) );
  INV3 U333 ( .A(A[22]), .Q(n172) );
  INV3 U334 ( .A(A[23]), .Q(n173) );
  CLKIN0 U335 ( .A(A[21]), .Q(n171) );
  INV3 U336 ( .A(A[26]), .Q(n176) );
  INV0 U337 ( .A(A[19]), .Q(n169) );
  INV0 U338 ( .A(A[30]), .Q(n180) );
  INV3 U339 ( .A(n149), .Q(n148) );
  NAND22 U340 ( .A(n150), .B(B[0]), .Q(n149) );
  INV0 U341 ( .A(A[0]), .Q(n150) );
  INV0 U342 ( .A(A[15]), .Q(n165) );
  INV0 U343 ( .A(A[24]), .Q(n174) );
  INV0 U344 ( .A(A[14]), .Q(n164) );
  INV0 U345 ( .A(A[11]), .Q(n161) );
  INV3 U346 ( .A(A[27]), .Q(n177) );
  INV0 U347 ( .A(A[17]), .Q(n167) );
  NAND22 U348 ( .A(B[13]), .B(n163), .Q(n87) );
  CLKIN0 U349 ( .A(A[18]), .Q(n168) );
  INV0 U350 ( .A(A[8]), .Q(n158) );
  NAND22 U351 ( .A(B[30]), .B(n180), .Q(n10) );
  CLKIN0 U352 ( .A(A[5]), .Q(n155) );
endmodule


module sqroot_seq_NBITS32_DW01_sub_5 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n45,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n62,
         n63, n64, n65, n66, n67, n68, n69, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n85, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n108, n109, n110, n111,
         n112, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n130, n131, n132, n133, n135, n137, n140, n141,
         n142, n143, n144, n146, n147, n148, n149, n150, n151, n152, n153,
         n156, n157, n158, n159, n160, n161, n162, n164, n165, n166, n167,
         n168, n169, n170, n171, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n195,
         n196, n197, n198, n199, n200, n203, n204, n205, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n220, n221,
         n222, n223, n224, n225, n227, n230, n231, n232, n233, n235, n236,
         n237, n238, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n258, n259, n260,
         n261, n262, n264, n265, n266, n268, n270, n271, n272, n273, n274,
         n275, n277, n278, n280, n283, n284, n285, n286, n287, n288, n289,
         n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459;

  OAI212 U22 ( .A(n48), .B(n83), .C(n49), .Q(n47) );
  OAI212 U26 ( .A(n62), .B(n52), .C(n53), .Q(n51) );
  OAI212 U32 ( .A(n55), .B(n459), .C(n56), .Q(n54) );
  OAI212 U36 ( .A(n59), .B(n69), .C(n62), .Q(n58) );
  OAI212 U44 ( .A(n64), .B(n459), .C(n65), .Q(n63) );
  OAI212 U52 ( .A(n80), .B(n72), .C(n73), .Q(n67) );
  OAI212 U58 ( .A(n75), .B(n459), .C(n76), .Q(n74) );
  OAI212 U68 ( .A(n82), .B(n459), .C(n83), .Q(n81) );
  AOI212 U74 ( .A(n103), .B(n88), .C(n89), .Q(n83) );
  OAI212 U76 ( .A(n98), .B(n90), .C(n91), .Q(n89) );
  OAI212 U82 ( .A(n93), .B(n459), .C(n94), .Q(n92) );
  OAI212 U92 ( .A(n100), .B(n459), .C(n101), .Q(n99) );
  OAI212 U100 ( .A(n112), .B(n108), .C(n109), .Q(n103) );
  OAI212 U114 ( .A(n151), .B(n116), .C(n117), .Q(n115) );
  AOI212 U116 ( .A(n135), .B(n118), .C(n119), .Q(n117) );
  OAI212 U118 ( .A(n130), .B(n120), .C(n121), .Q(n119) );
  OAI212 U144 ( .A(n148), .B(n140), .C(n141), .Q(n135) );
  OAI212 U150 ( .A(n143), .B(n430), .C(n144), .Q(n142) );
  AOI212 U166 ( .A(n156), .B(n171), .C(n157), .Q(n151) );
  OAI212 U174 ( .A(n161), .B(n430), .C(n162), .Q(n160) );
  OAI212 U192 ( .A(n180), .B(n176), .C(n177), .Q(n171) );
  NOR24 U195 ( .A(n309), .B(A[15]), .Q(n176) );
  AOI212 U207 ( .A(n185), .B(n198), .C(n186), .Q(n184) );
  OAI212 U209 ( .A(n195), .B(n187), .C(n188), .Q(n186) );
  NOR24 U212 ( .A(n311), .B(A[13]), .Q(n187) );
  XNR22 U244 ( .A(n25), .B(n216), .Q(DIFF[9]) );
  AOI212 U246 ( .A(n231), .B(n212), .C(n213), .Q(n211) );
  OAI212 U248 ( .A(n214), .B(n218), .C(n215), .Q(n213) );
  NOR24 U251 ( .A(n315), .B(A[9]), .Q(n214) );
  AOI212 U256 ( .A(n285), .B(n227), .C(n220), .Q(n218) );
  NOR24 U261 ( .A(n316), .B(A[8]), .Q(n221) );
  NOR24 U271 ( .A(n317), .B(A[7]), .Q(n224) );
  OAI212 U275 ( .A(n232), .B(n244), .C(n233), .Q(n231) );
  AOI212 U277 ( .A(n287), .B(n240), .C(n235), .Q(n233) );
  AOI212 U294 ( .A(n245), .B(n253), .C(n246), .Q(n244) );
  OAI212 U296 ( .A(n247), .B(n251), .C(n248), .Q(n246) );
  OAI212 U309 ( .A(n254), .B(n256), .C(n255), .Q(n253) );
  AOI212 U315 ( .A(n292), .B(n2), .C(n258), .Q(n256) );
  INV0 U360 ( .A(B[1]), .Q(n323) );
  OAI211 U361 ( .A(n250), .B(n252), .C(n251), .Q(n249) );
  NOR23 U362 ( .A(n214), .B(n217), .Q(n212) );
  BUF15 U363 ( .A(n1), .Q(n459) );
  INV0 U364 ( .A(n98), .Q(n96) );
  NAND21 U365 ( .A(n95), .B(n98), .Q(n10) );
  NAND23 U366 ( .A(A[24]), .B(n300), .Q(n98) );
  NOR22 U367 ( .A(n59), .B(n68), .Q(n57) );
  AOI212 U368 ( .A(n85), .B(n57), .C(n58), .Q(n56) );
  XNR22 U369 ( .A(n3), .B(n36), .Q(DIFF[31]) );
  INV6 U370 ( .A(n83), .Q(n85) );
  NOR23 U371 ( .A(n52), .B(n59), .Q(n50) );
  NOR22 U372 ( .A(n295), .B(A[29]), .Q(n52) );
  NAND24 U373 ( .A(n456), .B(n180), .Q(n178) );
  NOR22 U374 ( .A(n299), .B(A[25]), .Q(n90) );
  NOR23 U375 ( .A(n187), .B(n192), .Q(n185) );
  NAND22 U376 ( .A(n39), .B(n448), .Q(n449) );
  NOR22 U377 ( .A(n108), .B(n111), .Q(n102) );
  NAND22 U378 ( .A(A[12]), .B(n312), .Q(n195) );
  NOR21 U379 ( .A(n322), .B(A[2]), .Q(n254) );
  NAND22 U380 ( .A(A[3]), .B(n321), .Q(n251) );
  NAND22 U381 ( .A(A[8]), .B(n316), .Q(n222) );
  NAND22 U382 ( .A(n439), .B(n444), .Q(n149) );
  NAND22 U383 ( .A(n447), .B(n448), .Q(n451) );
  NAND22 U384 ( .A(A[5]), .B(n319), .Q(n242) );
  NAND23 U385 ( .A(A[18]), .B(n306), .Q(n148) );
  NAND23 U386 ( .A(A[20]), .B(n304), .Q(n130) );
  NAND21 U387 ( .A(n266), .B(n73), .Q(n7) );
  INV6 U388 ( .A(n183), .Q(n452) );
  BUF2 U389 ( .A(n187), .Q(n427) );
  NOR23 U390 ( .A(n300), .B(A[24]), .Q(n97) );
  NOR23 U391 ( .A(n320), .B(A[4]), .Q(n247) );
  NOR23 U392 ( .A(n310), .B(A[14]), .Q(n179) );
  CLKIN12 U393 ( .A(n181), .Q(n429) );
  NOR23 U394 ( .A(n140), .B(n147), .Q(n457) );
  NOR23 U395 ( .A(n306), .B(A[18]), .Q(n147) );
  NAND21 U396 ( .A(n77), .B(n80), .Q(n8) );
  CLKIN3 U397 ( .A(n80), .Q(n78) );
  CLKIN3 U398 ( .A(n457), .Q(n458) );
  NAND24 U399 ( .A(n457), .B(n118), .Q(n116) );
  NAND23 U400 ( .A(n287), .B(n288), .Q(n232) );
  INV3 U401 ( .A(n66), .Q(n68) );
  NAND22 U402 ( .A(A[25]), .B(n299), .Q(n91) );
  NAND24 U403 ( .A(n442), .B(n204), .Q(n198) );
  AOI211 U404 ( .A(n85), .B(n77), .C(n78), .Q(n76) );
  INV3 U405 ( .A(n449), .Q(n450) );
  NOR22 U406 ( .A(n296), .B(A[28]), .Q(n59) );
  INV3 U407 ( .A(n203), .Q(n441) );
  NAND22 U408 ( .A(A[22]), .B(n302), .Q(n112) );
  INV3 U409 ( .A(n48), .Q(n447) );
  INV3 U410 ( .A(n224), .Q(n286) );
  INV3 U411 ( .A(n222), .Q(n220) );
  INV3 U412 ( .A(n225), .Q(n227) );
  INV3 U413 ( .A(n241), .Q(n288) );
  NAND22 U414 ( .A(A[9]), .B(n315), .Q(n215) );
  XNR21 U415 ( .A(n26), .B(n223), .Q(DIFF[8]) );
  XOR20 U416 ( .A(n27), .B(n230), .Q(DIFF[7]) );
  INV6 U417 ( .A(n236), .Q(n287) );
  AOI211 U418 ( .A(n156), .B(n171), .C(n157), .Q(n428) );
  INV6 U419 ( .A(n211), .Q(n453) );
  NAND22 U420 ( .A(n102), .B(n88), .Q(n82) );
  INV3 U421 ( .A(n82), .Q(n448) );
  INV3 U422 ( .A(n166), .Q(n164) );
  INV1 U423 ( .A(n253), .Q(n252) );
  NAND28 U424 ( .A(n446), .B(n159), .Q(n157) );
  NOR24 U425 ( .A(n318), .B(A[6]), .Q(n236) );
  NAND22 U426 ( .A(n156), .B(n170), .Q(n150) );
  INV15 U427 ( .A(n429), .Q(n430) );
  NAND21 U428 ( .A(n297), .B(A[27]), .Q(n73) );
  AOI312 U429 ( .A(n431), .B(n432), .C(n182), .D(n115), .Q(n1) );
  INV6 U430 ( .A(n116), .Q(n431) );
  INV3 U431 ( .A(n150), .Q(n432) );
  NAND26 U432 ( .A(A[14]), .B(n310), .Q(n180) );
  NOR22 U433 ( .A(n176), .B(n179), .Q(n170) );
  INV1 U434 ( .A(n165), .Q(n277) );
  CLKIN6 U435 ( .A(n182), .Q(n181) );
  BUF2 U436 ( .A(n256), .Q(n433) );
  INV2 U437 ( .A(n192), .Q(n434) );
  INV3 U438 ( .A(n434), .Q(n435) );
  NOR23 U439 ( .A(n312), .B(A[12]), .Q(n192) );
  NAND21 U440 ( .A(n277), .B(n166), .Q(n18) );
  NAND21 U441 ( .A(n434), .B(n195), .Q(n22) );
  INV2 U442 ( .A(n428), .Q(n153) );
  NOR24 U443 ( .A(n79), .B(n72), .Q(n66) );
  NOR23 U444 ( .A(n298), .B(A[26]), .Q(n79) );
  AOI211 U445 ( .A(n85), .B(n66), .C(n67), .Q(n65) );
  INV0 U446 ( .A(n148), .Q(n146) );
  NAND26 U447 ( .A(n454), .B(n184), .Q(n182) );
  INV2 U448 ( .A(n231), .Q(n230) );
  CLKIN0 U449 ( .A(n127), .Q(n273) );
  OAI210 U450 ( .A(n435), .B(n200), .C(n195), .Q(n191) );
  NAND21 U451 ( .A(n275), .B(n148), .Q(n16) );
  NAND21 U452 ( .A(n152), .B(n457), .Q(n132) );
  BUF2 U453 ( .A(n445), .Q(n436) );
  NAND21 U454 ( .A(n280), .B(n188), .Q(n21) );
  BUF2 U455 ( .A(n225), .Q(n437) );
  NAND22 U456 ( .A(n152), .B(n438), .Q(n439) );
  INV2 U457 ( .A(n430), .Q(n438) );
  CLKIN1 U458 ( .A(n153), .Q(n444) );
  NAND21 U459 ( .A(A[19]), .B(n305), .Q(n141) );
  AOI212 U460 ( .A(n67), .B(n50), .C(n51), .Q(n49) );
  NAND22 U461 ( .A(A[11]), .B(n313), .Q(n204) );
  INV6 U462 ( .A(n209), .Q(n440) );
  INV0 U463 ( .A(n209), .Q(n207) );
  NAND26 U464 ( .A(A[10]), .B(n314), .Q(n209) );
  NAND22 U465 ( .A(A[21]), .B(n303), .Q(n121) );
  NOR24 U466 ( .A(n303), .B(A[21]), .Q(n120) );
  NAND24 U467 ( .A(n441), .B(n440), .Q(n442) );
  NAND24 U468 ( .A(n286), .B(n285), .Q(n217) );
  INV3 U469 ( .A(n200), .Q(n443) );
  CLKIN3 U470 ( .A(n198), .Q(n200) );
  NAND21 U471 ( .A(A[13]), .B(n311), .Q(n188) );
  NAND22 U472 ( .A(n448), .B(n57), .Q(n55) );
  NOR23 U473 ( .A(n203), .B(n208), .Q(n197) );
  NAND26 U474 ( .A(n453), .B(n452), .Q(n454) );
  INV1 U475 ( .A(n208), .Q(n283) );
  NOR23 U476 ( .A(n314), .B(A[10]), .Q(n208) );
  INV0 U477 ( .A(B[7]), .Q(n317) );
  NAND22 U478 ( .A(n125), .B(n152), .Q(n123) );
  INV2 U479 ( .A(n150), .Q(n152) );
  INV1 U480 ( .A(n147), .Q(n275) );
  NAND24 U481 ( .A(n164), .B(n445), .Q(n446) );
  CLKIN6 U482 ( .A(n158), .Q(n445) );
  NAND22 U483 ( .A(A[17]), .B(n307), .Q(n159) );
  XOR22 U484 ( .A(n21), .B(n189), .Q(DIFF[13]) );
  NOR20 U485 ( .A(n435), .B(n199), .Q(n190) );
  AOI212 U486 ( .A(n47), .B(n39), .C(n40), .Q(n38) );
  INV0 U487 ( .A(B[2]), .Q(n322) );
  CLKIN0 U488 ( .A(n176), .Q(n278) );
  NAND20 U489 ( .A(n278), .B(n177), .Q(n19) );
  NAND21 U490 ( .A(n455), .B(n180), .Q(n20) );
  NOR24 U491 ( .A(n297), .B(A[27]), .Q(n72) );
  NOR21 U492 ( .A(n127), .B(n458), .Q(n125) );
  INV4 U493 ( .A(n67), .Q(n69) );
  XOR21 U494 ( .A(n459), .B(n12), .Q(DIFF[22]) );
  AOI210 U495 ( .A(n153), .B(n457), .C(n135), .Q(n133) );
  NOR23 U496 ( .A(n321), .B(A[3]), .Q(n250) );
  NOR22 U497 ( .A(n250), .B(n247), .Q(n245) );
  XNR22 U498 ( .A(n17), .B(n160), .Q(DIFF[17]) );
  OAI211 U499 ( .A(n451), .B(n459), .C(n45), .Q(n43) );
  OAI211 U500 ( .A(n37), .B(n459), .C(n38), .Q(n36) );
  NAND24 U501 ( .A(n66), .B(n50), .Q(n48) );
  AOI212 U502 ( .A(n210), .B(n283), .C(n207), .Q(n205) );
  XOR22 U503 ( .A(n23), .B(n205), .Q(DIFF[11]) );
  NOR24 U504 ( .A(n127), .B(n120), .Q(n118) );
  XNR22 U505 ( .A(n8), .B(n81), .Q(DIFF[26]) );
  NAND21 U506 ( .A(A[15]), .B(n309), .Q(n177) );
  NAND24 U507 ( .A(n455), .B(n429), .Q(n456) );
  NAND21 U508 ( .A(n284), .B(n215), .Q(n25) );
  XNR22 U509 ( .A(n14), .B(n131), .Q(DIFF[20]) );
  OAI212 U510 ( .A(n132), .B(n430), .C(n133), .Q(n131) );
  XNR22 U511 ( .A(n6), .B(n63), .Q(DIFF[28]) );
  XNR22 U512 ( .A(n99), .B(n10), .Q(DIFF[24]) );
  XNR22 U513 ( .A(n15), .B(n142), .Q(DIFF[19]) );
  CLKIN2 U514 ( .A(n197), .Q(n199) );
  XNR22 U515 ( .A(n54), .B(n5), .Q(DIFF[29]) );
  NAND22 U516 ( .A(A[23]), .B(n301), .Q(n109) );
  NOR24 U517 ( .A(n313), .B(A[11]), .Q(n203) );
  CLKIN3 U518 ( .A(n259), .Q(n292) );
  XNR22 U519 ( .A(n13), .B(n122), .Q(DIFF[21]) );
  XNR22 U520 ( .A(n11), .B(n110), .Q(DIFF[23]) );
  OAI212 U521 ( .A(n217), .B(n230), .C(n218), .Q(n216) );
  XNR22 U522 ( .A(n9), .B(n92), .Q(DIFF[25]) );
  NOR24 U523 ( .A(n305), .B(A[19]), .Q(n140) );
  INV1 U524 ( .A(n135), .Q(n137) );
  OAI211 U525 ( .A(n127), .B(n137), .C(n130), .Q(n126) );
  INV4 U526 ( .A(n237), .Q(n235) );
  OAI211 U527 ( .A(n224), .B(n230), .C(n437), .Q(n223) );
  OAI212 U528 ( .A(n111), .B(n459), .C(n112), .Q(n110) );
  AOI211 U529 ( .A(n153), .B(n275), .C(n146), .Q(n144) );
  AOI211 U530 ( .A(n153), .B(n125), .C(n126), .Q(n124) );
  XNR22 U531 ( .A(n19), .B(n178), .Q(DIFF[15]) );
  NAND22 U532 ( .A(A[26]), .B(n298), .Q(n80) );
  AOI212 U533 ( .A(n243), .B(n288), .C(n240), .Q(n238) );
  INV1 U534 ( .A(n244), .Q(n243) );
  XOR22 U535 ( .A(n22), .B(n196), .Q(DIFF[12]) );
  AOI211 U536 ( .A(n210), .B(n197), .C(n443), .Q(n196) );
  XNR22 U537 ( .A(n7), .B(n74), .Q(DIFF[27]) );
  INV0 U538 ( .A(n111), .Q(n271) );
  NOR22 U539 ( .A(n302), .B(A[22]), .Q(n111) );
  XNR22 U540 ( .A(n18), .B(n167), .Q(DIFF[16]) );
  OAI212 U541 ( .A(n168), .B(n430), .C(n169), .Q(n167) );
  NOR22 U542 ( .A(n165), .B(n158), .Q(n156) );
  NOR24 U543 ( .A(n307), .B(A[17]), .Q(n158) );
  INV0 U544 ( .A(n214), .Q(n284) );
  AOI211 U545 ( .A(n210), .B(n190), .C(n191), .Q(n189) );
  XNR22 U546 ( .A(n16), .B(n149), .Q(DIFF[18]) );
  NOR22 U547 ( .A(n319), .B(A[5]), .Q(n241) );
  INV2 U548 ( .A(n211), .Q(n210) );
  INV3 U549 ( .A(n260), .Q(n258) );
  NAND23 U550 ( .A(A[6]), .B(n318), .Q(n237) );
  CLKIN3 U551 ( .A(n261), .Q(n2) );
  NAND22 U552 ( .A(n152), .B(n275), .Q(n143) );
  CLKIN0 U553 ( .A(n179), .Q(n455) );
  INV0 U554 ( .A(n120), .Q(n272) );
  CLKIN0 U555 ( .A(B[8]), .Q(n316) );
  XOR21 U556 ( .A(n20), .B(n430), .Q(DIFF[14]) );
  NAND24 U557 ( .A(n197), .B(n185), .Q(n183) );
  CLKIN0 U558 ( .A(n170), .Q(n168) );
  OAI212 U559 ( .A(n123), .B(n430), .C(n124), .Q(n122) );
  CLKIN1 U560 ( .A(n79), .Q(n77) );
  NAND20 U561 ( .A(n288), .B(n242), .Q(n29) );
  INV0 U562 ( .A(n72), .Q(n266) );
  INV0 U563 ( .A(n108), .Q(n270) );
  NAND21 U564 ( .A(A[31]), .B(n293), .Q(n35) );
  CLKIN0 U565 ( .A(B[0]), .Q(n324) );
  NAND21 U566 ( .A(n283), .B(n209), .Q(n24) );
  NAND22 U567 ( .A(n448), .B(n77), .Q(n75) );
  INV0 U568 ( .A(n140), .Q(n274) );
  INV0 U569 ( .A(n59), .Q(n265) );
  INV1 U570 ( .A(n97), .Q(n95) );
  NAND21 U571 ( .A(n39), .B(n42), .Q(n4) );
  INV0 U572 ( .A(n52), .Q(n264) );
  NOR24 U573 ( .A(n304), .B(A[20]), .Q(n127) );
  NAND21 U574 ( .A(A[28]), .B(n296), .Q(n62) );
  NOR21 U575 ( .A(n323), .B(A[1]), .Q(n259) );
  NAND21 U576 ( .A(A[30]), .B(n294), .Q(n42) );
  NAND20 U577 ( .A(A[29]), .B(n295), .Q(n53) );
  NAND22 U578 ( .A(A[2]), .B(n322), .Q(n255) );
  NAND21 U579 ( .A(A[1]), .B(n323), .Q(n260) );
  INV2 U580 ( .A(n34), .Q(n262) );
  CLKIN0 U581 ( .A(B[14]), .Q(n310) );
  CLKIN0 U582 ( .A(B[12]), .Q(n312) );
  CLKIN0 U583 ( .A(B[18]), .Q(n306) );
  CLKIN0 U584 ( .A(B[19]), .Q(n305) );
  XOR20 U585 ( .A(n261), .B(n33), .Q(DIFF[1]) );
  XNR20 U586 ( .A(n324), .B(A[0]), .Q(DIFF[0]) );
  INV0 U587 ( .A(B[27]), .Q(n297) );
  INV0 U588 ( .A(B[29]), .Q(n295) );
  INV0 U589 ( .A(n171), .Q(n169) );
  INV3 U590 ( .A(n102), .Q(n100) );
  INV0 U591 ( .A(n103), .Q(n101) );
  NAND22 U592 ( .A(n448), .B(n66), .Q(n64) );
  INV3 U593 ( .A(n47), .Q(n45) );
  NAND20 U594 ( .A(n287), .B(n237), .Q(n28) );
  NAND20 U595 ( .A(n170), .B(n277), .Q(n161) );
  AOI210 U596 ( .A(n171), .B(n277), .C(n164), .Q(n162) );
  NAND20 U597 ( .A(n102), .B(n95), .Q(n93) );
  AOI210 U598 ( .A(n103), .B(n95), .C(n96), .Q(n94) );
  NAND22 U599 ( .A(n262), .B(n35), .Q(n3) );
  NOR23 U600 ( .A(n90), .B(n97), .Q(n88) );
  INV3 U601 ( .A(n42), .Q(n40) );
  NAND20 U602 ( .A(n436), .B(n159), .Q(n17) );
  NAND20 U603 ( .A(n441), .B(n204), .Q(n23) );
  NAND22 U604 ( .A(n289), .B(n248), .Q(n30) );
  INV0 U605 ( .A(n247), .Q(n289) );
  NAND20 U606 ( .A(n273), .B(n130), .Q(n14) );
  NAND20 U607 ( .A(n274), .B(n141), .Q(n15) );
  INV3 U608 ( .A(n242), .Q(n240) );
  NAND20 U609 ( .A(n292), .B(n260), .Q(n33) );
  NAND20 U610 ( .A(n286), .B(n437), .Q(n27) );
  NAND22 U611 ( .A(n291), .B(n255), .Q(n32) );
  INV0 U612 ( .A(n254), .Q(n291) );
  NAND22 U613 ( .A(n265), .B(n62), .Q(n6) );
  NAND22 U614 ( .A(n264), .B(n53), .Q(n5) );
  NAND22 U615 ( .A(n272), .B(n121), .Q(n13) );
  NAND22 U616 ( .A(n270), .B(n109), .Q(n11) );
  NAND22 U617 ( .A(n268), .B(n91), .Q(n9) );
  INV0 U618 ( .A(n90), .Q(n268) );
  NAND22 U619 ( .A(n271), .B(n112), .Q(n12) );
  NAND22 U620 ( .A(n290), .B(n251), .Q(n31) );
  INV0 U621 ( .A(n250), .Q(n290) );
  INV0 U622 ( .A(n427), .Q(n280) );
  NAND22 U623 ( .A(n450), .B(n447), .Q(n37) );
  NAND22 U624 ( .A(A[4]), .B(n320), .Q(n248) );
  NOR23 U625 ( .A(n301), .B(A[23]), .Q(n108) );
  CLKIN0 U626 ( .A(B[6]), .Q(n318) );
  NAND24 U627 ( .A(A[7]), .B(n317), .Q(n225) );
  INV3 U628 ( .A(n41), .Q(n39) );
  NOR21 U629 ( .A(n294), .B(A[30]), .Q(n41) );
  NAND22 U630 ( .A(A[16]), .B(n308), .Q(n166) );
  NOR21 U631 ( .A(n324), .B(A[0]), .Q(n261) );
  NOR22 U632 ( .A(n308), .B(A[16]), .Q(n165) );
  NOR21 U633 ( .A(n293), .B(A[31]), .Q(n34) );
  CLKIN0 U634 ( .A(B[10]), .Q(n314) );
  CLKIN0 U635 ( .A(B[15]), .Q(n309) );
  XOR20 U636 ( .A(n433), .B(n32), .Q(DIFF[2]) );
  XNR21 U637 ( .A(n4), .B(n43), .Q(DIFF[30]) );
  XNR21 U638 ( .A(n29), .B(n243), .Q(DIFF[5]) );
  XNR21 U639 ( .A(n30), .B(n249), .Q(DIFF[4]) );
  CLKIN0 U640 ( .A(B[3]), .Q(n321) );
  XOR21 U641 ( .A(n28), .B(n238), .Q(DIFF[6]) );
  XOR21 U642 ( .A(n31), .B(n252), .Q(DIFF[3]) );
  XNR21 U643 ( .A(n24), .B(n210), .Q(DIFF[10]) );
  INV0 U644 ( .A(B[22]), .Q(n302) );
  CLKIN0 U645 ( .A(B[16]), .Q(n308) );
  INV0 U646 ( .A(B[28]), .Q(n296) );
  INV0 U647 ( .A(B[26]), .Q(n298) );
  INV0 U648 ( .A(B[21]), .Q(n303) );
  INV0 U649 ( .A(B[25]), .Q(n299) );
  INV0 U650 ( .A(B[24]), .Q(n300) );
  CLKIN0 U651 ( .A(B[13]), .Q(n311) );
  INV0 U652 ( .A(B[23]), .Q(n301) );
  INV0 U653 ( .A(B[20]), .Q(n304) );
  INV0 U654 ( .A(B[17]), .Q(n307) );
  INV3 U655 ( .A(B[31]), .Q(n293) );
  INV3 U656 ( .A(B[30]), .Q(n294) );
  INV0 U657 ( .A(B[9]), .Q(n315) );
  CLKIN0 U658 ( .A(B[4]), .Q(n320) );
  INV0 U659 ( .A(B[11]), .Q(n313) );
  INV1 U660 ( .A(B[5]), .Q(n319) );
  NAND20 U661 ( .A(n285), .B(n222), .Q(n26) );
  CLKIN6 U662 ( .A(n221), .Q(n285) );
endmodule


module sqroot_seq_NBITS32_DW_cmp_6 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, 
        EQ_NE );
  input [31:0] A;
  input [31:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n249, n250,
         n251;

  OAI212 U1 ( .A(n1), .B(n25), .C(n2), .Q(GE_LT_GT_LE) );
  AOI212 U3 ( .A(n8), .B(n3), .C(n4), .Q(n2) );
  OAI212 U9 ( .A(n9), .B(n12), .C(n10), .Q(n8) );
  AOI212 U13 ( .A(n20), .B(n13), .C(n14), .Q(n12) );
  OAI212 U15 ( .A(n18), .B(n15), .C(n16), .Q(n14) );
  OAI212 U21 ( .A(n21), .B(n24), .C(n22), .Q(n20) );
  AOI212 U26 ( .A(n56), .B(n26), .C(n27), .Q(n25) );
  OAI212 U28 ( .A(n28), .B(n43), .C(n29), .Q(n27) );
  OAI212 U32 ( .A(n35), .B(n32), .C(n33), .Q(n31) );
  NOR24 U33 ( .A(B[25]), .B(n169), .Q(n32) );
  OAI212 U38 ( .A(n41), .B(n38), .C(n39), .Q(n37) );
  OAI212 U46 ( .A(n49), .B(n46), .C(n47), .Q(n45) );
  OAI212 U52 ( .A(n55), .B(n52), .C(n53), .Q(n51) );
  OAI212 U57 ( .A(n57), .B(n87), .C(n58), .Q(n56) );
  OAI212 U61 ( .A(n64), .B(n61), .C(n62), .Q(n60) );
  OAI212 U67 ( .A(n78), .B(n67), .C(n68), .Q(n66) );
  AOI212 U79 ( .A(n79), .B(n84), .C(n80), .Q(n78) );
  AOI212 U88 ( .A(n110), .B(n88), .C(n89), .Q(n87) );
  OAI212 U90 ( .A(n101), .B(n90), .C(n91), .Q(n89) );
  AOI212 U102 ( .A(n102), .B(n107), .C(n103), .Q(n101) );
  OAI212 U111 ( .A(n111), .B(n121), .C(n112), .Q(n110) );
  OAI212 U124 ( .A(n127), .B(n124), .C(n125), .Q(n123) );
  OAI212 U129 ( .A(n129), .B(n131), .C(n130), .Q(n128) );
  OAI212 U137 ( .A(n139), .B(n137), .C(n138), .Q(n136) );
  INV3 U180 ( .A(n82), .Q(n80) );
  INV8 U181 ( .A(A[23]), .Q(n167) );
  NOR23 U182 ( .A(B[23]), .B(n167), .Q(n38) );
  INV3 U183 ( .A(A[11]), .Q(n155) );
  NAND23 U184 ( .A(n170), .B(B[26]), .Q(n24) );
  INV3 U185 ( .A(A[21]), .Q(n165) );
  NOR22 U186 ( .A(n149), .B(B[5]), .Q(n124) );
  INV6 U187 ( .A(A[27]), .Q(n171) );
  NAND23 U188 ( .A(B[24]), .B(n168), .Q(n35) );
  INV3 U189 ( .A(n105), .Q(n103) );
  AOI211 U190 ( .A(n92), .B(n97), .C(n93), .Q(n91) );
  NOR22 U191 ( .A(n157), .B(B[13]), .Q(n81) );
  NOR23 U192 ( .A(B[27]), .B(n171), .Q(n21) );
  CLKIN3 U193 ( .A(A[26]), .Q(n170) );
  NOR23 U194 ( .A(B[19]), .B(n163), .Q(n52) );
  NOR22 U195 ( .A(B[31]), .B(n175), .Q(n5) );
  INV3 U196 ( .A(A[9]), .Q(n153) );
  NAND23 U197 ( .A(n96), .B(n92), .Q(n90) );
  NOR24 U198 ( .A(n250), .B(n40), .Q(n36) );
  CLKIN12 U199 ( .A(A[29]), .Q(n173) );
  INV3 U200 ( .A(n95), .Q(n93) );
  NOR22 U201 ( .A(n9), .B(n11), .Q(n7) );
  INV3 U202 ( .A(A[20]), .Q(n164) );
  NOR22 U203 ( .A(n63), .B(n61), .Q(n59) );
  INV3 U204 ( .A(A[31]), .Q(n175) );
  NAND21 U205 ( .A(n175), .B(B[31]), .Q(n6) );
  NOR23 U206 ( .A(n159), .B(B[15]), .Q(n71) );
  AOI212 U207 ( .A(n44), .B(n51), .C(n45), .Q(n43) );
  NOR22 U208 ( .A(n77), .B(n67), .Q(n65) );
  NAND24 U209 ( .A(n69), .B(n73), .Q(n67) );
  NAND24 U210 ( .A(n166), .B(B[22]), .Q(n41) );
  NOR23 U211 ( .A(n46), .B(n48), .Q(n44) );
  NOR24 U212 ( .A(B[21]), .B(n165), .Q(n46) );
  NAND22 U213 ( .A(n164), .B(B[20]), .Q(n49) );
  NOR24 U214 ( .A(B[30]), .B(n174), .Q(n9) );
  NOR23 U215 ( .A(B[9]), .B(n153), .Q(n104) );
  CLKIN6 U216 ( .A(n94), .Q(n92) );
  NAND21 U217 ( .A(n174), .B(B[30]), .Q(n10) );
  NOR23 U218 ( .A(n42), .B(n28), .Q(n26) );
  NAND21 U219 ( .A(n165), .B(B[21]), .Q(n47) );
  NOR21 U220 ( .A(B[27]), .B(n171), .Q(n249) );
  NOR23 U221 ( .A(B[28]), .B(n172), .Q(n17) );
  NOR24 U222 ( .A(n34), .B(n251), .Q(n30) );
  CLKIN6 U223 ( .A(A[17]), .Q(n161) );
  CLKIN4 U224 ( .A(A[30]), .Q(n174) );
  NAND21 U225 ( .A(n163), .B(B[19]), .Q(n53) );
  NOR22 U226 ( .A(B[26]), .B(n170), .Q(n23) );
  CLKIN6 U227 ( .A(A[14]), .Q(n158) );
  NAND21 U228 ( .A(n161), .B(B[17]), .Q(n62) );
  AOI212 U229 ( .A(n30), .B(n37), .C(n31), .Q(n29) );
  NOR22 U230 ( .A(B[23]), .B(n167), .Q(n250) );
  AOI212 U231 ( .A(n128), .B(n122), .C(n123), .Q(n121) );
  CLKIN6 U232 ( .A(A[22]), .Q(n166) );
  NOR23 U233 ( .A(B[14]), .B(n158), .Q(n75) );
  NOR23 U234 ( .A(B[22]), .B(n166), .Q(n40) );
  NOR23 U235 ( .A(n17), .B(n15), .Q(n13) );
  NOR23 U236 ( .A(n169), .B(B[25]), .Q(n251) );
  CLKIN12 U237 ( .A(A[25]), .Q(n169) );
  NAND23 U238 ( .A(n19), .B(n13), .Q(n11) );
  NAND24 U239 ( .A(n36), .B(n30), .Q(n28) );
  NOR24 U240 ( .A(n168), .B(B[24]), .Q(n34) );
  NAND22 U241 ( .A(n162), .B(B[18]), .Q(n55) );
  AOI212 U242 ( .A(n69), .B(n74), .C(n70), .Q(n68) );
  NOR22 U243 ( .A(B[12]), .B(n156), .Q(n85) );
  NAND23 U244 ( .A(n156), .B(B[12]), .Q(n86) );
  NOR21 U245 ( .A(n52), .B(n54), .Q(n50) );
  NAND22 U246 ( .A(B[15]), .B(n159), .Q(n72) );
  INV6 U247 ( .A(n75), .Q(n73) );
  NAND21 U248 ( .A(n171), .B(B[27]), .Q(n22) );
  NOR22 U249 ( .A(n23), .B(n249), .Q(n19) );
  CLKIN6 U250 ( .A(n71), .Q(n69) );
  CLKIN6 U251 ( .A(A[15]), .Q(n159) );
  NAND21 U252 ( .A(n153), .B(B[9]), .Q(n105) );
  NOR24 U253 ( .A(B[17]), .B(n161), .Q(n61) );
  NOR23 U254 ( .A(B[11]), .B(n155), .Q(n94) );
  NAND22 U255 ( .A(n158), .B(B[14]), .Q(n76) );
  NOR24 U256 ( .A(B[29]), .B(n173), .Q(n15) );
  NOR22 U257 ( .A(B[18]), .B(n162), .Q(n54) );
  NAND21 U258 ( .A(n144), .B(B[0]), .Q(n143) );
  CLKIN2 U259 ( .A(n142), .Q(n140) );
  CLKIN2 U260 ( .A(n116), .Q(n114) );
  CLKIN3 U261 ( .A(n72), .Q(n70) );
  CLKIN2 U262 ( .A(A[1]), .Q(n145) );
  NAND21 U263 ( .A(n146), .B(B[2]), .Q(n135) );
  CLKIN3 U264 ( .A(A[12]), .Q(n156) );
  CLKIN3 U265 ( .A(A[6]), .Q(n150) );
  AOI212 U266 ( .A(n66), .B(n59), .C(n60), .Q(n58) );
  NAND22 U267 ( .A(n83), .B(n79), .Q(n77) );
  CLKIN3 U268 ( .A(n85), .Q(n83) );
  INV3 U269 ( .A(n5), .Q(n3) );
  CLKIN3 U270 ( .A(A[8]), .Q(n152) );
  CLKIN3 U271 ( .A(A[10]), .Q(n154) );
  CLKIN3 U272 ( .A(A[5]), .Q(n149) );
  INV2 U273 ( .A(n6), .Q(n4) );
  CLKIN2 U274 ( .A(A[4]), .Q(n148) );
  CLKIN3 U275 ( .A(n134), .Q(n132) );
  CLKIN3 U276 ( .A(A[7]), .Q(n151) );
  CLKIN3 U277 ( .A(A[2]), .Q(n146) );
  CLKIN3 U278 ( .A(A[3]), .Q(n147) );
  NAND20 U279 ( .A(n151), .B(B[7]), .Q(n116) );
  NAND21 U280 ( .A(n154), .B(B[10]), .Q(n99) );
  NAND21 U281 ( .A(n152), .B(B[8]), .Q(n109) );
  NAND21 U282 ( .A(n150), .B(B[6]), .Q(n120) );
  NOR20 U283 ( .A(B[0]), .B(n144), .Q(n142) );
  NAND21 U284 ( .A(n148), .B(B[4]), .Q(n127) );
  NAND20 U285 ( .A(n147), .B(B[3]), .Q(n130) );
  NAND20 U286 ( .A(n145), .B(B[1]), .Q(n138) );
  CLKIN3 U287 ( .A(n115), .Q(n113) );
  CLKIN3 U288 ( .A(A[13]), .Q(n157) );
  NOR21 U289 ( .A(n126), .B(n124), .Q(n122) );
  NOR21 U290 ( .A(n100), .B(n90), .Q(n88) );
  AOI211 U291 ( .A(n136), .B(n132), .C(n133), .Q(n131) );
  INV3 U292 ( .A(n135), .Q(n133) );
  INV3 U293 ( .A(A[19]), .Q(n163) );
  CLKIN3 U294 ( .A(A[16]), .Q(n160) );
  INV3 U295 ( .A(A[0]), .Q(n144) );
  NAND22 U296 ( .A(n65), .B(n59), .Q(n57) );
  CLKIN3 U297 ( .A(A[18]), .Q(n162) );
  NAND22 U298 ( .A(n7), .B(n3), .Q(n1) );
  NOR21 U299 ( .A(B[4]), .B(n148), .Q(n126) );
  NOR21 U300 ( .A(B[2]), .B(n146), .Q(n134) );
  NOR21 U301 ( .A(B[7]), .B(n151), .Q(n115) );
  NOR22 U302 ( .A(n160), .B(B[16]), .Q(n63) );
  NOR21 U303 ( .A(B[1]), .B(n145), .Q(n137) );
  NOR21 U304 ( .A(B[3]), .B(n147), .Q(n129) );
  CLKIN3 U305 ( .A(n109), .Q(n107) );
  CLKIN3 U306 ( .A(n76), .Q(n74) );
  CLKIN3 U307 ( .A(n99), .Q(n97) );
  AOI211 U308 ( .A(n113), .B(n118), .C(n114), .Q(n112) );
  CLKIN3 U309 ( .A(n120), .Q(n118) );
  NAND20 U310 ( .A(n149), .B(B[5]), .Q(n125) );
  CLKIN3 U311 ( .A(n104), .Q(n102) );
  CLKIN3 U312 ( .A(n98), .Q(n96) );
  NOR21 U313 ( .A(B[10]), .B(n154), .Q(n98) );
  NAND21 U314 ( .A(n102), .B(n106), .Q(n100) );
  CLKIN3 U315 ( .A(n108), .Q(n106) );
  NOR21 U316 ( .A(B[8]), .B(n152), .Q(n108) );
  NAND22 U317 ( .A(n50), .B(n44), .Q(n42) );
  NOR21 U318 ( .A(n141), .B(n140), .Q(n139) );
  INV3 U319 ( .A(n143), .Q(n141) );
  NAND22 U320 ( .A(n113), .B(n117), .Q(n111) );
  CLKIN3 U321 ( .A(n119), .Q(n117) );
  NOR21 U322 ( .A(B[6]), .B(n150), .Q(n119) );
  CLKIN3 U323 ( .A(n86), .Q(n84) );
  NAND22 U324 ( .A(B[16]), .B(n160), .Q(n64) );
  NAND21 U325 ( .A(n157), .B(B[13]), .Q(n82) );
  NAND21 U326 ( .A(n155), .B(B[11]), .Q(n95) );
  NAND21 U327 ( .A(n173), .B(B[29]), .Q(n16) );
  NAND21 U328 ( .A(n167), .B(B[23]), .Q(n39) );
  NAND22 U329 ( .A(n172), .B(B[28]), .Q(n18) );
  NAND21 U330 ( .A(B[25]), .B(n169), .Q(n33) );
  NOR22 U331 ( .A(B[20]), .B(n164), .Q(n48) );
  CLKIN6 U332 ( .A(n81), .Q(n79) );
  CLKIN6 U333 ( .A(A[28]), .Q(n172) );
  CLKIN6 U334 ( .A(A[24]), .Q(n168) );
endmodule


module sqroot_seq_NBITS32_DW01_add_5 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n50, n51, n52, n54, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n67, n68, n69, n70, n73, n74, n75, n76, n77, n78, n79,
         n80, n83, n84, n85, n86, n87, n88, n90, n91, n92, n93, n94, n96, n99,
         n100, n101, n102, n103, n104, n105, n107, n108, n109, n110, n111,
         n112, n113, n114, n119, n120, n121, n122, n123, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n141, n142, n143, n144, n145, n146, n147, n148, n151, n152, n153,
         n154, n155, n158, n159, n160, n161, n162, n163, n164, n167, n168,
         n169, n170, n171, n172, n173, n175, n176, n177, n178, n179, n180,
         n181, n182, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n206, n207, n208,
         n209, n210, n211, n214, n215, n216, n217, n218, n219, n220, n222,
         n223, n224, n225, n227, n228, n229, n230, n231, n232, n233, n234,
         n235, n237, n239, n240, n241, n242, n246, n247, n248, n249, n250,
         n251, n252, n253, n257, n258, n259, n260, n261, n262, n264, n267,
         n268, n269, n270, n272, n273, n274, n275, n277, n278, n279, n280,
         n281, n283, n284, n285, n286, n287, n288, n291, n292, n295, n297,
         n298, n299, n300, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n313, n314, n315, n316, n317, n318, n319, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479;

  XNR22 U30 ( .A(n4), .B(n65), .Q(SUM[28]) );
  OAI212 U35 ( .A(n59), .B(n94), .C(n60), .Q(n58) );
  AOI212 U47 ( .A(n96), .B(n68), .C(n69), .Q(n67) );
  OAI212 U49 ( .A(n70), .B(n80), .C(n73), .Q(n69) );
  OAI212 U57 ( .A(n75), .B(n479), .C(n76), .Q(n74) );
  AOI212 U87 ( .A(n114), .B(n99), .C(n100), .Q(n94) );
  OAI212 U89 ( .A(n109), .B(n101), .C(n102), .Q(n100) );
  OAI212 U95 ( .A(n104), .B(n479), .C(n105), .Q(n103) );
  OAI212 U113 ( .A(n123), .B(n119), .C(n120), .Q(n114) );
  OAI212 U119 ( .A(n122), .B(n479), .C(n123), .Q(n121) );
  AOI212 U125 ( .A(n125), .B(n193), .C(n126), .Q(n1) );
  OAI212 U127 ( .A(n162), .B(n127), .C(n128), .Q(n126) );
  AOI212 U129 ( .A(n146), .B(n129), .C(n130), .Q(n128) );
  OAI212 U131 ( .A(n131), .B(n141), .C(n132), .Q(n130) );
  NOR24 U146 ( .A(B[19]), .B(A[19]), .Q(n138) );
  AOI212 U179 ( .A(n182), .B(n167), .C(n168), .Q(n162) );
  OAI212 U181 ( .A(n177), .B(n169), .C(n170), .Q(n168) );
  NOR24 U194 ( .A(B[15]), .B(A[15]), .Q(n176) );
  OAI212 U197 ( .A(n192), .B(n179), .C(n180), .Q(n178) );
  OAI212 U205 ( .A(n191), .B(n187), .C(n188), .Q(n182) );
  NOR24 U208 ( .A(B[14]), .B(A[14]), .Q(n187) );
  OAI212 U211 ( .A(n192), .B(n190), .C(n191), .Q(n189) );
  AOI212 U220 ( .A(n209), .B(n196), .C(n197), .Q(n195) );
  OAI212 U222 ( .A(n206), .B(n198), .C(n199), .Q(n197) );
  NOR24 U235 ( .A(B[11]), .B(A[11]), .Q(n203) );
  OAI212 U244 ( .A(n214), .B(n220), .C(n215), .Q(n209) );
  AOI212 U254 ( .A(n310), .B(n227), .C(n222), .Q(n220) );
  AOI212 U271 ( .A(n268), .B(n232), .C(n233), .Q(n231) );
  OAI212 U273 ( .A(n251), .B(n234), .C(n235), .Q(n233) );
  OAI212 U320 ( .A(n281), .B(n269), .C(n270), .Q(n268) );
  AOI212 U322 ( .A(n316), .B(n277), .C(n272), .Q(n270) );
  CLKIN6 U355 ( .A(n50), .Q(n3) );
  CLKIN6 U356 ( .A(n42), .Q(n40) );
  AOI211 U357 ( .A(n58), .B(n50), .C(n51), .Q(n47) );
  CLKIN6 U358 ( .A(A[29]), .Q(n52) );
  OAI211 U359 ( .A(n203), .B(n211), .C(n206), .Q(n202) );
  NOR24 U360 ( .A(n158), .B(n422), .Q(n145) );
  NOR23 U361 ( .A(A[2]), .B(B[2]), .Q(n278) );
  INV6 U362 ( .A(n262), .Q(n264) );
  CLKIN4 U363 ( .A(n284), .Q(n318) );
  NAND28 U364 ( .A(n470), .B(n152), .Q(n146) );
  NAND24 U365 ( .A(n181), .B(n167), .Q(n161) );
  NOR23 U366 ( .A(B[18]), .B(A[18]), .Q(n422) );
  NOR24 U367 ( .A(B[21]), .B(A[21]), .Q(n122) );
  NAND26 U368 ( .A(n56), .B(n478), .Q(n54) );
  CLKIN8 U369 ( .A(n247), .Q(n313) );
  NAND21 U370 ( .A(n74), .B(n5), .Q(n429) );
  INV4 U371 ( .A(n74), .Q(n428) );
  CLKIN6 U372 ( .A(n258), .Q(n314) );
  NOR23 U373 ( .A(n452), .B(n108), .Q(n99) );
  NOR23 U374 ( .A(B[23]), .B(A[23]), .Q(n108) );
  NOR23 U375 ( .A(B[17]), .B(A[17]), .Q(n158) );
  CLKIN6 U376 ( .A(n223), .Q(n310) );
  NAND24 U377 ( .A(A[17]), .B(B[17]), .Q(n159) );
  NOR22 U378 ( .A(B[25]), .B(A[25]), .Q(n90) );
  INV3 U379 ( .A(n5), .Q(n427) );
  NAND26 U380 ( .A(A[21]), .B(B[21]), .Q(n123) );
  AOI211 U381 ( .A(n78), .B(n61), .C(n62), .Q(n60) );
  INV3 U382 ( .A(n248), .Q(n246) );
  INV3 U383 ( .A(n229), .Q(n227) );
  NOR23 U384 ( .A(B[10]), .B(A[10]), .Q(n214) );
  INV3 U385 ( .A(n77), .Q(n79) );
  NOR23 U386 ( .A(B[22]), .B(A[22]), .Q(n119) );
  NOR23 U387 ( .A(B[13]), .B(A[13]), .Q(n190) );
  NAND24 U388 ( .A(A[13]), .B(B[13]), .Q(n191) );
  NAND22 U389 ( .A(n77), .B(n61), .Q(n59) );
  NOR22 U390 ( .A(n451), .B(n461), .Q(n144) );
  NOR23 U391 ( .A(n450), .B(n147), .Q(n451) );
  NAND22 U392 ( .A(n424), .B(n438), .Q(n426) );
  INV3 U393 ( .A(n52), .Q(n50) );
  NAND23 U394 ( .A(n429), .B(n430), .Q(SUM[27]) );
  XNR21 U395 ( .A(n33), .B(n34), .Q(SUM[31]) );
  NOR24 U396 ( .A(B[20]), .B(A[20]), .Q(n131) );
  NAND22 U397 ( .A(B[7]), .B(A[7]), .Q(n239) );
  INV1 U398 ( .A(n114), .Q(n112) );
  NAND28 U399 ( .A(n475), .B(n112), .Q(n110) );
  NAND26 U400 ( .A(n469), .B(n468), .Q(n470) );
  NAND23 U401 ( .A(n311), .B(n310), .Q(n219) );
  NOR23 U402 ( .A(n214), .B(n219), .Q(n208) );
  AOI212 U403 ( .A(n96), .B(n88), .C(n431), .Q(n87) );
  NOR23 U404 ( .A(n234), .B(n250), .Q(n232) );
  NOR22 U405 ( .A(n93), .B(n463), .Q(n462) );
  INV1 U406 ( .A(n147), .Q(n423) );
  NAND22 U407 ( .A(n178), .B(n17), .Q(n425) );
  NAND22 U408 ( .A(n425), .B(n426), .Q(SUM[15]) );
  INV3 U409 ( .A(n178), .Q(n424) );
  NAND24 U410 ( .A(n427), .B(n428), .Q(n430) );
  NAND22 U411 ( .A(n292), .B(n73), .Q(n5) );
  INV3 U412 ( .A(n162), .Q(n164) );
  XOR22 U413 ( .A(n23), .B(n225), .Q(SUM[9]) );
  AOI212 U414 ( .A(n230), .B(n208), .C(n439), .Q(n207) );
  NAND23 U415 ( .A(n208), .B(n196), .Q(n194) );
  CLKIN6 U416 ( .A(n92), .Q(n465) );
  NAND26 U417 ( .A(n477), .B(n437), .Q(n92) );
  XOR22 U418 ( .A(n11), .B(n479), .Q(SUM[21]) );
  INV6 U419 ( .A(n54), .Q(n454) );
  NAND26 U420 ( .A(n455), .B(n456), .Q(SUM[29]) );
  INV0 U421 ( .A(n220), .Q(n218) );
  NAND24 U422 ( .A(A[11]), .B(B[11]), .Q(n206) );
  AOI210 U423 ( .A(n164), .B(n302), .C(n468), .Q(n155) );
  INV6 U424 ( .A(n164), .Q(n450) );
  INV6 U425 ( .A(n193), .Q(n192) );
  NAND22 U426 ( .A(n57), .B(n37), .Q(n35) );
  NAND24 U427 ( .A(n57), .B(n474), .Q(n478) );
  NOR22 U428 ( .A(n59), .B(n93), .Q(n57) );
  INV1 U429 ( .A(n113), .Q(n111) );
  NAND23 U430 ( .A(n113), .B(n99), .Q(n93) );
  NOR23 U431 ( .A(n119), .B(n122), .Q(n113) );
  NAND22 U432 ( .A(B[9]), .B(A[9]), .Q(n224) );
  NOR22 U433 ( .A(n70), .B(n79), .Q(n68) );
  AOI211 U434 ( .A(n58), .B(n37), .C(n38), .Q(n36) );
  INV3 U435 ( .A(n228), .Q(n311) );
  XOR21 U436 ( .A(n28), .B(n267), .Q(SUM[4]) );
  INV3 U437 ( .A(n250), .Q(n252) );
  INV3 U438 ( .A(B[7]), .Q(n460) );
  NOR22 U439 ( .A(n63), .B(n70), .Q(n61) );
  NAND22 U440 ( .A(n431), .B(n432), .Q(n433) );
  INV3 U441 ( .A(n70), .Q(n292) );
  INV3 U442 ( .A(n68), .Q(n463) );
  INV3 U443 ( .A(n17), .Q(n438) );
  CLKIN6 U444 ( .A(n110), .Q(n441) );
  INV3 U445 ( .A(n9), .Q(n440) );
  NAND22 U446 ( .A(n434), .B(n444), .Q(n436) );
  NAND23 U447 ( .A(A[19]), .B(B[19]), .Q(n141) );
  NAND22 U448 ( .A(n476), .B(n88), .Q(n86) );
  INV2 U449 ( .A(n474), .Q(n449) );
  NAND26 U450 ( .A(n454), .B(n453), .Q(n456) );
  NAND26 U451 ( .A(n313), .B(n458), .Q(n234) );
  NOR22 U452 ( .A(n138), .B(n147), .Q(n136) );
  NAND22 U453 ( .A(A[18]), .B(B[18]), .Q(n152) );
  INV6 U454 ( .A(n159), .Q(n468) );
  NAND26 U455 ( .A(n433), .B(n84), .Q(n78) );
  CLKIN3 U456 ( .A(n91), .Q(n431) );
  CLKIN3 U457 ( .A(n83), .Q(n432) );
  NAND22 U458 ( .A(n103), .B(n8), .Q(n435) );
  NAND22 U459 ( .A(n435), .B(n436), .Q(SUM[24]) );
  INV3 U460 ( .A(n103), .Q(n434) );
  CLKIN1 U461 ( .A(n209), .Q(n211) );
  XOR31 U462 ( .A(A[30]), .B(B[30]), .C(n45), .Q(SUM[30]) );
  NAND24 U463 ( .A(n474), .B(n462), .Q(n472) );
  XNR21 U464 ( .A(n14), .B(n153), .Q(SUM[18]) );
  XNR21 U465 ( .A(n16), .B(n171), .Q(SUM[16]) );
  INV2 U466 ( .A(n96), .Q(n437) );
  OAI212 U467 ( .A(n35), .B(n449), .C(n36), .Q(n34) );
  INV6 U468 ( .A(A[7]), .Q(n459) );
  INV2 U469 ( .A(n211), .Q(n439) );
  INV3 U470 ( .A(n39), .Q(n37) );
  NAND23 U471 ( .A(A[23]), .B(B[23]), .Q(n109) );
  INV3 U472 ( .A(n8), .Q(n444) );
  NAND22 U473 ( .A(n9), .B(n110), .Q(n442) );
  NAND24 U474 ( .A(n440), .B(n441), .Q(n443) );
  NAND24 U475 ( .A(n442), .B(n443), .Q(SUM[23]) );
  OAI212 U476 ( .A(n46), .B(n449), .C(n47), .Q(n45) );
  NAND21 U477 ( .A(n57), .B(n50), .Q(n46) );
  NAND24 U478 ( .A(B[4]), .B(A[4]), .Q(n262) );
  INV0 U479 ( .A(n251), .Q(n253) );
  NAND24 U480 ( .A(n448), .B(n445), .Q(n446) );
  NAND21 U481 ( .A(n15), .B(n160), .Q(n447) );
  NAND24 U482 ( .A(n446), .B(n447), .Q(SUM[17]) );
  INV3 U483 ( .A(n160), .Q(n445) );
  INV3 U484 ( .A(n15), .Q(n448) );
  INV2 U485 ( .A(n161), .Q(n163) );
  CLKIN6 U486 ( .A(n151), .Q(n469) );
  OAI212 U487 ( .A(n172), .B(n192), .C(n173), .Q(n171) );
  AOI212 U488 ( .A(n96), .B(n77), .C(n78), .Q(n76) );
  INV3 U489 ( .A(n94), .Q(n96) );
  NAND26 U490 ( .A(n472), .B(n67), .Q(n65) );
  INV15 U491 ( .A(n479), .Q(n474) );
  NAND23 U492 ( .A(n315), .B(n314), .Q(n250) );
  NOR23 U493 ( .A(A[6]), .B(B[6]), .Q(n247) );
  INV3 U494 ( .A(n78), .Q(n80) );
  INV2 U495 ( .A(n63), .Q(n291) );
  NOR24 U496 ( .A(B[28]), .B(A[28]), .Q(n63) );
  NOR22 U497 ( .A(n161), .B(n127), .Q(n125) );
  NOR23 U498 ( .A(A[5]), .B(B[5]), .Q(n258) );
  NAND21 U499 ( .A(n423), .B(n163), .Q(n143) );
  INV1 U500 ( .A(n158), .Q(n302) );
  NAND22 U501 ( .A(n300), .B(n141), .Q(n13) );
  XNR22 U502 ( .A(n13), .B(n142), .Q(SUM[19]) );
  INV1 U503 ( .A(n148), .Q(n461) );
  OAI212 U504 ( .A(n154), .B(n192), .C(n155), .Q(n153) );
  NAND24 U505 ( .A(n129), .B(n145), .Q(n127) );
  NOR24 U506 ( .A(B[24]), .B(A[24]), .Q(n452) );
  NAND22 U507 ( .A(A[24]), .B(B[24]), .Q(n102) );
  NAND23 U508 ( .A(n474), .B(n476), .Q(n477) );
  NAND23 U509 ( .A(n317), .B(n316), .Q(n269) );
  NAND22 U510 ( .A(B[2]), .B(A[2]), .Q(n279) );
  NAND22 U511 ( .A(n54), .B(n3), .Q(n455) );
  INV3 U512 ( .A(n3), .Q(n453) );
  INV2 U513 ( .A(n180), .Q(n457) );
  INV1 U514 ( .A(n182), .Q(n180) );
  NAND21 U515 ( .A(A[14]), .B(B[14]), .Q(n188) );
  INV2 U516 ( .A(n145), .Q(n147) );
  NAND28 U517 ( .A(n459), .B(n460), .Q(n458) );
  INV3 U518 ( .A(n259), .Q(n257) );
  NAND28 U519 ( .A(A[15]), .B(B[15]), .Q(n177) );
  NOR24 U520 ( .A(n131), .B(n138), .Q(n129) );
  NAND21 U521 ( .A(A[16]), .B(B[16]), .Q(n170) );
  NAND21 U522 ( .A(n295), .B(n102), .Q(n8) );
  INV0 U523 ( .A(n198), .Q(n307) );
  NAND26 U524 ( .A(n466), .B(n467), .Q(SUM[25]) );
  NOR24 U525 ( .A(B[26]), .B(A[26]), .Q(n83) );
  OAI212 U526 ( .A(n73), .B(n63), .C(n64), .Q(n62) );
  NOR24 U527 ( .A(B[24]), .B(A[24]), .Q(n101) );
  XNR22 U528 ( .A(n6), .B(n85), .Q(SUM[26]) );
  NAND26 U529 ( .A(n474), .B(n473), .Q(n475) );
  INV1 U530 ( .A(n176), .Q(n304) );
  XNR22 U531 ( .A(n18), .B(n189), .Q(SUM[14]) );
  NOR24 U532 ( .A(A[9]), .B(B[9]), .Q(n223) );
  OAI210 U533 ( .A(n250), .B(n267), .C(n251), .Q(n249) );
  INV2 U534 ( .A(n146), .Q(n148) );
  INV2 U535 ( .A(n58), .Q(n56) );
  NAND22 U536 ( .A(A[12]), .B(B[12]), .Q(n199) );
  OAI212 U537 ( .A(n86), .B(n479), .C(n87), .Q(n85) );
  INV0 U538 ( .A(n131), .Q(n299) );
  NOR24 U539 ( .A(A[3]), .B(B[3]), .Q(n273) );
  XOR22 U540 ( .A(n21), .B(n207), .Q(SUM[11]) );
  INV3 U541 ( .A(n231), .Q(n230) );
  INV3 U542 ( .A(n93), .Q(n476) );
  XOR22 U543 ( .A(n20), .B(n200), .Q(SUM[12]) );
  AOI212 U544 ( .A(n230), .B(n201), .C(n202), .Q(n200) );
  NOR21 U545 ( .A(n203), .B(n210), .Q(n201) );
  NAND22 U546 ( .A(A[22]), .B(B[22]), .Q(n120) );
  NAND22 U547 ( .A(A[27]), .B(B[27]), .Q(n73) );
  NAND22 U548 ( .A(A[28]), .B(B[28]), .Q(n64) );
  NAND22 U549 ( .A(B[3]), .B(A[3]), .Q(n274) );
  NAND22 U550 ( .A(n7), .B(n92), .Q(n466) );
  NAND24 U551 ( .A(n465), .B(n464), .Q(n467) );
  INV3 U552 ( .A(n7), .Q(n464) );
  NAND20 U553 ( .A(n88), .B(n91), .Q(n7) );
  NAND21 U554 ( .A(A[26]), .B(B[26]), .Q(n84) );
  NOR24 U555 ( .A(n169), .B(n176), .Q(n167) );
  OAI212 U556 ( .A(n194), .B(n231), .C(n195), .Q(n193) );
  AOI211 U557 ( .A(n136), .B(n164), .C(n137), .Q(n135) );
  AOI212 U558 ( .A(n230), .B(n311), .C(n227), .Q(n225) );
  OAI211 U559 ( .A(n138), .B(n148), .C(n141), .Q(n137) );
  NAND22 U560 ( .A(A[25]), .B(B[25]), .Q(n91) );
  OAI211 U561 ( .A(n261), .B(n267), .C(n262), .Q(n260) );
  OAI211 U562 ( .A(n241), .B(n267), .C(n242), .Q(n240) );
  INV3 U563 ( .A(n268), .Q(n267) );
  NAND20 U564 ( .A(n291), .B(n64), .Q(n4) );
  NOR24 U565 ( .A(B[27]), .B(A[27]), .Q(n70) );
  NAND21 U566 ( .A(n302), .B(n159), .Q(n15) );
  NAND22 U567 ( .A(n476), .B(n77), .Q(n75) );
  NOR24 U568 ( .A(n83), .B(n90), .Q(n77) );
  CLKIN2 U569 ( .A(n108), .Q(n471) );
  NOR24 U570 ( .A(n198), .B(n203), .Q(n196) );
  INV2 U571 ( .A(n111), .Q(n473) );
  BUF15 U572 ( .A(n1), .Q(n479) );
  NOR22 U573 ( .A(A[8]), .B(B[8]), .Q(n228) );
  INV0 U574 ( .A(n119), .Q(n297) );
  NAND22 U575 ( .A(A[10]), .B(B[10]), .Q(n215) );
  AOI212 U576 ( .A(n314), .B(n264), .C(n257), .Q(n251) );
  NAND22 U577 ( .A(n163), .B(n302), .Q(n154) );
  NAND20 U578 ( .A(n432), .B(n84), .Q(n6) );
  NOR21 U579 ( .A(B[30]), .B(A[30]), .Q(n43) );
  AOI212 U580 ( .A(n230), .B(n217), .C(n218), .Q(n216) );
  XNR21 U581 ( .A(n24), .B(n230), .Q(SUM[8]) );
  CLKIN0 U582 ( .A(n181), .Q(n179) );
  AOI212 U583 ( .A(n318), .B(n286), .C(n283), .Q(n281) );
  CLKIN3 U584 ( .A(n285), .Q(n283) );
  AOI212 U585 ( .A(n246), .B(n458), .C(n237), .Q(n235) );
  CLKIN6 U586 ( .A(n239), .Q(n237) );
  XNR22 U587 ( .A(n10), .B(n121), .Q(SUM[22]) );
  NAND20 U588 ( .A(n305), .B(n188), .Q(n18) );
  CLKIN3 U589 ( .A(n261), .Q(n315) );
  NAND20 U590 ( .A(n314), .B(n259), .Q(n27) );
  INV0 U591 ( .A(n109), .Q(n107) );
  INV0 U592 ( .A(n452), .Q(n295) );
  CLKIN0 U593 ( .A(n177), .Q(n175) );
  INV0 U594 ( .A(n138), .Q(n300) );
  NAND20 U595 ( .A(n471), .B(n109), .Q(n9) );
  NAND20 U596 ( .A(n458), .B(n239), .Q(n25) );
  XNR20 U597 ( .A(n286), .B(n31), .Q(SUM[1]) );
  NAND20 U598 ( .A(n318), .B(n285), .Q(n31) );
  NOR24 U599 ( .A(B[12]), .B(A[12]), .Q(n198) );
  NOR24 U600 ( .A(B[18]), .B(A[18]), .Q(n151) );
  NOR24 U601 ( .A(B[16]), .B(A[16]), .Q(n169) );
  NOR22 U602 ( .A(A[1]), .B(B[1]), .Q(n284) );
  NAND22 U603 ( .A(B[0]), .B(A[0]), .Q(n288) );
  NAND22 U604 ( .A(A[30]), .B(B[30]), .Q(n44) );
  NOR20 U605 ( .A(A[0]), .B(B[0]), .Q(n287) );
  NAND22 U606 ( .A(n113), .B(n471), .Q(n104) );
  NAND22 U607 ( .A(n136), .B(n163), .Q(n134) );
  NAND20 U608 ( .A(n181), .B(n304), .Q(n172) );
  INV3 U609 ( .A(n219), .Q(n217) );
  NAND20 U610 ( .A(n306), .B(n191), .Q(n19) );
  INV0 U611 ( .A(n190), .Q(n306) );
  INV3 U612 ( .A(n274), .Q(n272) );
  INV3 U613 ( .A(n224), .Q(n222) );
  NAND22 U614 ( .A(n297), .B(n120), .Q(n10) );
  NAND22 U615 ( .A(n307), .B(n199), .Q(n20) );
  NAND20 U616 ( .A(n298), .B(n123), .Q(n11) );
  INV3 U617 ( .A(n122), .Q(n298) );
  INV3 U618 ( .A(n90), .Q(n88) );
  XNR21 U619 ( .A(n25), .B(n240), .Q(SUM[7]) );
  NAND20 U620 ( .A(n311), .B(n229), .Q(n24) );
  AOI210 U621 ( .A(n114), .B(n471), .C(n107), .Q(n105) );
  AOI210 U622 ( .A(n457), .B(n304), .C(n175), .Q(n173) );
  NAND20 U623 ( .A(n252), .B(n313), .Q(n241) );
  XNR21 U624 ( .A(n26), .B(n249), .Q(SUM[6]) );
  NAND20 U625 ( .A(n313), .B(n248), .Q(n26) );
  XNR21 U626 ( .A(n30), .B(n280), .Q(SUM[2]) );
  NAND20 U627 ( .A(n317), .B(n279), .Q(n30) );
  XNR21 U628 ( .A(n27), .B(n260), .Q(SUM[5]) );
  NAND20 U629 ( .A(n310), .B(n224), .Q(n23) );
  XOR21 U630 ( .A(n29), .B(n275), .Q(SUM[3]) );
  NAND20 U631 ( .A(n316), .B(n274), .Q(n29) );
  AOI210 U632 ( .A(n280), .B(n317), .C(n277), .Q(n275) );
  XOR21 U633 ( .A(n22), .B(n216), .Q(SUM[10]) );
  NAND22 U634 ( .A(n309), .B(n215), .Q(n22) );
  NAND20 U635 ( .A(n315), .B(n262), .Q(n28) );
  INV3 U636 ( .A(n169), .Q(n303) );
  CLKIN0 U637 ( .A(n208), .Q(n210) );
  XNR21 U638 ( .A(n12), .B(n133), .Q(SUM[20]) );
  NAND20 U639 ( .A(n299), .B(n132), .Q(n12) );
  INV3 U640 ( .A(n288), .Q(n286) );
  INV0 U641 ( .A(n203), .Q(n308) );
  NAND22 U642 ( .A(n303), .B(n170), .Q(n16) );
  INV3 U643 ( .A(n279), .Q(n277) );
  INV0 U644 ( .A(n214), .Q(n309) );
  INV3 U645 ( .A(n32), .Q(SUM[0]) );
  NAND22 U646 ( .A(n319), .B(n288), .Q(n32) );
  INV3 U647 ( .A(n287), .Q(n319) );
  NAND22 U648 ( .A(n308), .B(n206), .Q(n21) );
  NAND22 U649 ( .A(n304), .B(n177), .Q(n17) );
  NAND22 U650 ( .A(B[5]), .B(A[5]), .Q(n259) );
  NOR23 U651 ( .A(A[4]), .B(B[4]), .Q(n261) );
  INV3 U652 ( .A(n43), .Q(n41) );
  NAND22 U653 ( .A(B[1]), .B(A[1]), .Q(n285) );
  NAND22 U654 ( .A(A[6]), .B(B[6]), .Q(n248) );
  INV3 U655 ( .A(A[31]), .Q(n33) );
  NAND22 U656 ( .A(n50), .B(n41), .Q(n39) );
  CLKIN3 U657 ( .A(n40), .Q(n38) );
  CLKIN3 U658 ( .A(n44), .Q(n42) );
  LOGIC0 U659 ( .Q(n51) );
  OAI211 U660 ( .A(n161), .B(n192), .C(n450), .Q(n160) );
  NAND20 U661 ( .A(n152), .B(n469), .Q(n14) );
  INV2 U662 ( .A(n187), .Q(n305) );
  NOR22 U663 ( .A(n187), .B(n190), .Q(n181) );
  AOI210 U664 ( .A(n253), .B(n313), .C(n246), .Q(n242) );
  INV2 U665 ( .A(n281), .Q(n280) );
  NAND24 U666 ( .A(B[8]), .B(A[8]), .Q(n229) );
  NAND22 U667 ( .A(A[20]), .B(B[20]), .Q(n132) );
  OAI212 U668 ( .A(n134), .B(n192), .C(n135), .Q(n133) );
  OAI212 U669 ( .A(n143), .B(n192), .C(n144), .Q(n142) );
  XOR21 U670 ( .A(n192), .B(n19), .Q(SUM[13]) );
  CLKIN6 U671 ( .A(n278), .Q(n317) );
  CLKIN6 U672 ( .A(n273), .Q(n316) );
endmodule


module sqroot_seq_NBITS32_DW01_add_6 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n68, n69, n70, n71, n72, n73, n74, n75,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n106, n107,
         n108, n109, n110, n111, n112, n113, n116, n117, n118, n119, n120,
         n122, n123, n124, n125, n126, n127, n128, n129, n132, n133, n134,
         n135, n136, n137, n138, n140, n141, n142, n143, n144, n145, n146,
         n147, n152, n153, n154, n155, n156, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n174, n175,
         n176, n177, n178, n179, n180, n181, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n200, n201, n202,
         n203, n204, n205, n206, n208, n209, n210, n211, n212, n213, n214,
         n215, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n239, n240, n241, n242,
         n243, n244, n247, n248, n249, n251, n252, n253, n254, n255, n256,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n269, n271, n272, n273, n274, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n425;

  OAI212 U22 ( .A(n47), .B(n55), .C(n48), .Q(n46) );
  XNR22 U27 ( .A(n7), .B(n60), .Q(SUM[28]) );
  AOI212 U34 ( .A(n73), .B(n56), .C(n57), .Q(n55) );
  OAI212 U36 ( .A(n68), .B(n58), .C(n59), .Q(n57) );
  OAI212 U42 ( .A(n61), .B(n415), .C(n62), .Q(n60) );
  XNR22 U53 ( .A(n9), .B(n80), .Q(SUM[26]) );
  OAI212 U62 ( .A(n86), .B(n78), .C(n79), .Q(n73) );
  XNR22 U77 ( .A(n11), .B(n98), .Q(SUM[24]) );
  OAI212 U82 ( .A(n92), .B(n127), .C(n93), .Q(n2) );
  OAI212 U86 ( .A(n106), .B(n96), .C(n97), .Q(n95) );
  XNR22 U91 ( .A(n12), .B(n107), .Q(SUM[23]) );
  XNR22 U103 ( .A(n13), .B(n118), .Q(SUM[22]) );
  OAI212 U112 ( .A(n124), .B(n116), .C(n117), .Q(n111) );
  XNR22 U117 ( .A(n14), .B(n125), .Q(SUM[21]) );
  OAI212 U118 ( .A(n119), .B(n425), .C(n120), .Q(n118) );
  XNR22 U127 ( .A(n136), .B(n15), .Q(SUM[20]) );
  AOI212 U134 ( .A(n147), .B(n132), .C(n133), .Q(n127) );
  OAI212 U136 ( .A(n142), .B(n134), .C(n135), .Q(n133) );
  XNR22 U141 ( .A(n16), .B(n143), .Q(SUM[19]) );
  OAI212 U142 ( .A(n137), .B(n425), .C(n138), .Q(n136) );
  XNR22 U151 ( .A(n154), .B(n17), .Q(SUM[18]) );
  OAI212 U152 ( .A(n144), .B(n425), .C(n145), .Q(n143) );
  OAI212 U160 ( .A(n156), .B(n152), .C(n153), .Q(n147) );
  OAI212 U166 ( .A(n155), .B(n425), .C(n156), .Q(n154) );
  XNR22 U171 ( .A(n166), .B(n19), .Q(SUM[16]) );
  OAI212 U174 ( .A(n195), .B(n160), .C(n161), .Q(n159) );
  AOI212 U176 ( .A(n179), .B(n162), .C(n163), .Q(n161) );
  XNR22 U183 ( .A(n20), .B(n175), .Q(SUM[15]) );
  NOR24 U193 ( .A(B[15]), .B(A[15]), .Q(n171) );
  XNR22 U195 ( .A(n21), .B(n186), .Q(SUM[14]) );
  OAI212 U204 ( .A(n192), .B(n184), .C(n185), .Q(n179) );
  OAI212 U210 ( .A(n187), .B(n225), .C(n188), .Q(n186) );
  AOI212 U226 ( .A(n215), .B(n200), .C(n201), .Q(n195) );
  OAI212 U228 ( .A(n210), .B(n202), .C(n203), .Q(n201) );
  OAI212 U244 ( .A(n212), .B(n225), .C(n213), .Q(n211) );
  OAI212 U252 ( .A(n224), .B(n220), .C(n221), .Q(n215) );
  OAI212 U258 ( .A(n223), .B(n225), .C(n224), .Q(n222) );
  OAI212 U265 ( .A(n255), .B(n227), .C(n228), .Q(n226) );
  AOI212 U267 ( .A(n242), .B(n229), .C(n230), .Q(n228) );
  OAI212 U269 ( .A(n239), .B(n231), .C(n232), .Q(n230) );
  OAI212 U277 ( .A(n236), .B(n244), .C(n239), .Q(n235) );
  NOR24 U282 ( .A(B[7]), .B(A[7]), .Q(n236) );
  OAI212 U291 ( .A(n247), .B(n253), .C(n248), .Q(n242) );
  AOI212 U306 ( .A(n404), .B(n256), .C(n257), .Q(n255) );
  CLKIN6 U334 ( .A(n38), .Q(n5) );
  CLKIN6 U335 ( .A(A[30]), .Q(n40) );
  AOI210 U336 ( .A(n42), .B(n38), .C(n39), .Q(n37) );
  NOR22 U337 ( .A(B[19]), .B(A[19]), .Q(n141) );
  INV3 U338 ( .A(n264), .Q(n263) );
  NAND23 U339 ( .A(n403), .B(n416), .Q(n193) );
  NOR24 U340 ( .A(n171), .B(n164), .Q(n162) );
  NOR23 U341 ( .A(n261), .B(n258), .Q(n256) );
  OAI211 U342 ( .A(n65), .B(n75), .C(n68), .Q(n64) );
  NOR22 U343 ( .A(n65), .B(n58), .Q(n56) );
  OAI211 U344 ( .A(n50), .B(n415), .C(n51), .Q(n49) );
  NOR23 U345 ( .A(n422), .B(n64), .Q(n62) );
  NOR23 U346 ( .A(n134), .B(n141), .Q(n132) );
  OAI212 U347 ( .A(n81), .B(n425), .C(n82), .Q(n80) );
  OAI212 U348 ( .A(n99), .B(n425), .C(n100), .Q(n98) );
  CLKIN4 U349 ( .A(n2), .Q(n89) );
  AOI211 U350 ( .A(n2), .B(n83), .C(n84), .Q(n82) );
  XNR22 U351 ( .A(n5), .B(n42), .Q(SUM[30]) );
  AOI211 U352 ( .A(n129), .B(n101), .C(n102), .Q(n100) );
  NAND21 U353 ( .A(n3), .B(n83), .Q(n81) );
  NOR24 U354 ( .A(n92), .B(n126), .Q(n3) );
  INV2 U355 ( .A(n126), .Q(n128) );
  NAND24 U356 ( .A(n146), .B(n132), .Q(n126) );
  NAND22 U357 ( .A(A[5]), .B(B[5]), .Q(n253) );
  NOR23 U358 ( .A(n202), .B(n209), .Q(n200) );
  NOR21 U359 ( .A(n96), .B(n103), .Q(n94) );
  NAND23 U360 ( .A(n408), .B(n177), .Q(n175) );
  NOR21 U361 ( .A(B[26]), .B(A[26]), .Q(n78) );
  NOR21 U362 ( .A(B[27]), .B(A[27]), .Q(n65) );
  NOR21 U363 ( .A(B[28]), .B(A[28]), .Q(n58) );
  NOR21 U364 ( .A(n47), .B(n54), .Q(n45) );
  XNR21 U365 ( .A(n24), .B(n211), .Q(SUM[11]) );
  NAND21 U366 ( .A(A[25]), .B(B[25]), .Q(n86) );
  INV6 U367 ( .A(n225), .Q(n407) );
  BUF2 U368 ( .A(n266), .Q(n401) );
  NOR23 U369 ( .A(n423), .B(n78), .Q(n72) );
  OAI211 U370 ( .A(n108), .B(n425), .C(n109), .Q(n107) );
  CLKIN6 U371 ( .A(n241), .Q(n243) );
  INV3 U372 ( .A(n127), .Q(n129) );
  AOI211 U373 ( .A(n129), .B(n110), .C(n111), .Q(n109) );
  XNR21 U374 ( .A(n10), .B(n87), .Q(SUM[25]) );
  OAI212 U375 ( .A(n88), .B(n425), .C(n89), .Q(n87) );
  NAND22 U376 ( .A(n402), .B(n407), .Q(n403) );
  INV3 U377 ( .A(n194), .Q(n402) );
  NAND24 U378 ( .A(n214), .B(n200), .Q(n194) );
  CLKIN1 U379 ( .A(n197), .Q(n416) );
  NOR23 U380 ( .A(B[4]), .B(A[4]), .Q(n258) );
  NAND22 U381 ( .A(B[4]), .B(A[4]), .Q(n259) );
  XOR22 U382 ( .A(n18), .B(n425), .Q(SUM[17]) );
  NAND21 U383 ( .A(n3), .B(n45), .Q(n43) );
  NOR23 U384 ( .A(B[13]), .B(A[13]), .Q(n191) );
  INV3 U385 ( .A(n26), .Q(n413) );
  NAND22 U386 ( .A(A[21]), .B(B[21]), .Q(n124) );
  NOR23 U387 ( .A(B[11]), .B(A[11]), .Q(n209) );
  INV3 U388 ( .A(n194), .Q(n196) );
  INV3 U389 ( .A(n178), .Q(n180) );
  NOR22 U390 ( .A(B[18]), .B(A[18]), .Q(n152) );
  NOR22 U391 ( .A(B[17]), .B(A[17]), .Q(n155) );
  NAND22 U392 ( .A(A[17]), .B(B[17]), .Q(n156) );
  NAND22 U393 ( .A(A[19]), .B(B[19]), .Q(n142) );
  BUF2 U394 ( .A(n85), .Q(n423) );
  NOR23 U395 ( .A(n236), .B(n231), .Q(n229) );
  NOR21 U396 ( .A(n65), .B(n74), .Q(n63) );
  INV3 U397 ( .A(n72), .Q(n74) );
  AOI211 U398 ( .A(n111), .B(n94), .C(n95), .Q(n93) );
  INV3 U399 ( .A(n29), .Q(n412) );
  NAND22 U400 ( .A(A[11]), .B(B[11]), .Q(n210) );
  NAND22 U401 ( .A(n410), .B(n206), .Q(n204) );
  NOR23 U402 ( .A(B[14]), .B(A[14]), .Q(n184) );
  NOR23 U403 ( .A(B[22]), .B(A[22]), .Q(n116) );
  AOI211 U404 ( .A(n129), .B(n279), .C(n122), .Q(n120) );
  NOR22 U405 ( .A(B[23]), .B(A[23]), .Q(n103) );
  NOR22 U406 ( .A(B[24]), .B(A[24]), .Q(n96) );
  INV2 U407 ( .A(n34), .Q(SUM[1]) );
  NAND22 U408 ( .A(n298), .B(n401), .Q(n33) );
  NAND24 U409 ( .A(B[2]), .B(A[2]), .Q(n266) );
  INV3 U410 ( .A(n255), .Q(n254) );
  OAI211 U411 ( .A(n268), .B(n265), .C(n266), .Q(n264) );
  XNR21 U412 ( .A(n8), .B(n69), .Q(SUM[27]) );
  NAND21 U413 ( .A(n290), .B(n221), .Q(n25) );
  OAI212 U414 ( .A(n268), .B(n265), .C(n266), .Q(n404) );
  BUF2 U415 ( .A(n258), .Q(n405) );
  INV1 U416 ( .A(n242), .Q(n244) );
  NOR24 U417 ( .A(B[6]), .B(A[6]), .Q(n247) );
  CLKIN3 U418 ( .A(n425), .Q(n414) );
  INV6 U419 ( .A(n414), .Q(n415) );
  CLKIN3 U420 ( .A(n405), .Q(n296) );
  NAND24 U421 ( .A(n406), .B(n407), .Q(n408) );
  INV3 U422 ( .A(n176), .Q(n406) );
  NAND24 U423 ( .A(A[1]), .B(B[1]), .Q(n268) );
  NAND22 U424 ( .A(n407), .B(n409), .Q(n410) );
  INV3 U425 ( .A(n205), .Q(n409) );
  NOR22 U426 ( .A(B[10]), .B(A[10]), .Q(n220) );
  NOR24 U427 ( .A(B[12]), .B(A[12]), .Q(n202) );
  BUF2 U428 ( .A(n248), .Q(n411) );
  OAI210 U429 ( .A(n224), .B(n220), .C(n221), .Q(n418) );
  NOR23 U430 ( .A(n223), .B(n220), .Q(n214) );
  XNR22 U431 ( .A(n249), .B(n412), .Q(SUM[6]) );
  XNR22 U432 ( .A(n413), .B(n225), .Q(SUM[9]) );
  AOI212 U433 ( .A(n197), .B(n169), .C(n170), .Q(n168) );
  XNR22 U434 ( .A(n25), .B(n222), .Q(SUM[10]) );
  NOR23 U435 ( .A(B[9]), .B(A[9]), .Q(n223) );
  NAND21 U436 ( .A(n294), .B(n411), .Q(n29) );
  CLKIN0 U437 ( .A(n220), .Q(n290) );
  NAND21 U438 ( .A(n297), .B(n262), .Q(n32) );
  NOR24 U439 ( .A(n419), .B(n243), .Q(n420) );
  INV2 U440 ( .A(n179), .Q(n181) );
  NOR24 U441 ( .A(n420), .B(n417), .Q(n240) );
  NAND22 U442 ( .A(A[14]), .B(B[14]), .Q(n185) );
  NAND21 U443 ( .A(A[24]), .B(B[24]), .Q(n97) );
  CLKIN6 U444 ( .A(n254), .Q(n419) );
  XNR22 U445 ( .A(n23), .B(n204), .Q(SUM[12]) );
  CLKIN8 U446 ( .A(n226), .Q(n225) );
  XOR22 U447 ( .A(n27), .B(n233), .Q(SUM[8]) );
  INV0 U448 ( .A(n265), .Q(n298) );
  BUF2 U449 ( .A(n242), .Q(n417) );
  NOR24 U450 ( .A(A[2]), .B(B[2]), .Q(n265) );
  NAND21 U451 ( .A(A[20]), .B(B[20]), .Q(n135) );
  NAND23 U452 ( .A(A[9]), .B(B[9]), .Q(n224) );
  NAND21 U453 ( .A(A[16]), .B(B[16]), .Q(n165) );
  NOR24 U454 ( .A(B[16]), .B(A[16]), .Q(n164) );
  OAI210 U455 ( .A(n103), .B(n113), .C(n106), .Q(n102) );
  INV0 U456 ( .A(n103), .Q(n277) );
  OAI212 U457 ( .A(n167), .B(n225), .C(n168), .Q(n166) );
  NAND21 U458 ( .A(n3), .B(n72), .Q(n70) );
  XNR21 U459 ( .A(n31), .B(n260), .Q(SUM[4]) );
  AOI212 U460 ( .A(n254), .B(n295), .C(n251), .Q(n249) );
  INV3 U461 ( .A(n252), .Q(n295) );
  OAI211 U462 ( .A(n171), .B(n181), .C(n174), .Q(n170) );
  OAI212 U463 ( .A(n174), .B(n164), .C(n165), .Q(n163) );
  NAND22 U464 ( .A(A[15]), .B(B[15]), .Q(n174) );
  AOI210 U465 ( .A(n418), .B(n289), .C(n208), .Q(n206) );
  CLKIN0 U466 ( .A(n418), .Q(n213) );
  NAND21 U467 ( .A(n128), .B(n101), .Q(n99) );
  NAND22 U468 ( .A(n128), .B(n279), .Q(n119) );
  NAND22 U469 ( .A(n128), .B(n110), .Q(n108) );
  NAND21 U470 ( .A(n284), .B(n165), .Q(n19) );
  AOI212 U471 ( .A(n197), .B(n287), .C(n190), .Q(n188) );
  AOI211 U472 ( .A(n197), .B(n178), .C(n179), .Q(n177) );
  INV2 U473 ( .A(n195), .Q(n197) );
  XNR22 U474 ( .A(n22), .B(n193), .Q(SUM[13]) );
  NAND21 U475 ( .A(A[10]), .B(B[10]), .Q(n221) );
  NAND22 U476 ( .A(A[13]), .B(B[13]), .Q(n192) );
  INV2 U477 ( .A(n123), .Q(n279) );
  NOR22 U478 ( .A(B[21]), .B(A[21]), .Q(n123) );
  NOR24 U479 ( .A(n191), .B(n184), .Q(n178) );
  XOR21 U480 ( .A(n32), .B(n263), .Q(SUM[3]) );
  NAND20 U481 ( .A(n282), .B(n153), .Q(n17) );
  NAND21 U482 ( .A(A[18]), .B(B[18]), .Q(n153) );
  NAND21 U483 ( .A(A[6]), .B(B[6]), .Q(n248) );
  OAI211 U484 ( .A(n126), .B(n425), .C(n127), .Q(n125) );
  CLKBU15 U485 ( .A(n1), .Q(n425) );
  NOR23 U486 ( .A(n252), .B(n247), .Q(n241) );
  XOR22 U487 ( .A(n28), .B(n240), .Q(SUM[7]) );
  OAI211 U488 ( .A(n261), .B(n263), .C(n262), .Q(n260) );
  NAND22 U489 ( .A(A[3]), .B(B[3]), .Q(n262) );
  NOR24 U490 ( .A(n89), .B(n421), .Q(n422) );
  CLKIN3 U491 ( .A(n63), .Q(n421) );
  NAND21 U492 ( .A(A[12]), .B(B[12]), .Q(n203) );
  NOR21 U493 ( .A(n103), .B(n112), .Q(n101) );
  NAND20 U494 ( .A(n3), .B(n52), .Q(n50) );
  NAND21 U495 ( .A(n196), .B(n178), .Q(n176) );
  NAND21 U496 ( .A(n3), .B(n63), .Q(n61) );
  INV0 U497 ( .A(n236), .Q(n293) );
  OAI212 U498 ( .A(n262), .B(n258), .C(n259), .Q(n257) );
  INV3 U499 ( .A(n54), .Q(n52) );
  INV3 U500 ( .A(n55), .Q(n53) );
  CLKIN3 U501 ( .A(n73), .Q(n75) );
  CLKIN0 U502 ( .A(n65), .Q(n273) );
  NAND20 U503 ( .A(n273), .B(n68), .Q(n8) );
  CLKIN2 U504 ( .A(n3), .Q(n88) );
  NAND20 U505 ( .A(n83), .B(n86), .Q(n10) );
  CLKIN0 U506 ( .A(n111), .Q(n113) );
  NAND20 U507 ( .A(n280), .B(n135), .Q(n15) );
  INV0 U508 ( .A(n47), .Q(n271) );
  NAND21 U509 ( .A(n271), .B(n48), .Q(n6) );
  NAND21 U510 ( .A(A[23]), .B(B[23]), .Q(n106) );
  NAND21 U511 ( .A(A[22]), .B(B[22]), .Q(n117) );
  XNR21 U512 ( .A(n30), .B(n254), .Q(SUM[5]) );
  AOI212 U513 ( .A(n254), .B(n234), .C(n235), .Q(n233) );
  NAND21 U514 ( .A(n196), .B(n287), .Q(n187) );
  NAND20 U515 ( .A(n146), .B(n281), .Q(n137) );
  CLKIN0 U516 ( .A(n146), .Q(n144) );
  NOR20 U517 ( .A(n236), .B(n243), .Q(n234) );
  NOR21 U518 ( .A(n171), .B(n180), .Q(n169) );
  INV0 U519 ( .A(n134), .Q(n280) );
  CLKIN0 U520 ( .A(n110), .Q(n112) );
  INV0 U521 ( .A(n261), .Q(n297) );
  INV0 U522 ( .A(n96), .Q(n276) );
  NAND21 U523 ( .A(n287), .B(n192), .Q(n22) );
  NAND21 U524 ( .A(A[8]), .B(B[8]), .Q(n232) );
  NOR20 U525 ( .A(B[25]), .B(A[25]), .Q(n85) );
  NAND20 U526 ( .A(A[27]), .B(B[27]), .Q(n68) );
  NAND20 U527 ( .A(A[26]), .B(B[26]), .Q(n79) );
  NAND20 U528 ( .A(A[28]), .B(B[28]), .Q(n59) );
  NAND20 U529 ( .A(A[29]), .B(B[29]), .Q(n48) );
  NAND22 U530 ( .A(n72), .B(n56), .Q(n54) );
  NAND22 U531 ( .A(n110), .B(n94), .Q(n92) );
  NAND22 U532 ( .A(n196), .B(n169), .Q(n167) );
  NAND20 U533 ( .A(n214), .B(n289), .Q(n205) );
  CLKIN0 U534 ( .A(n214), .Q(n212) );
  NOR23 U535 ( .A(n123), .B(n116), .Q(n110) );
  NAND22 U536 ( .A(n241), .B(n229), .Q(n227) );
  NOR22 U537 ( .A(n152), .B(n155), .Q(n146) );
  NAND20 U538 ( .A(n283), .B(n156), .Q(n18) );
  INV3 U539 ( .A(n155), .Q(n283) );
  NAND20 U540 ( .A(n293), .B(n239), .Q(n28) );
  INV0 U541 ( .A(n247), .Q(n294) );
  INV0 U542 ( .A(n210), .Q(n208) );
  INV3 U543 ( .A(n423), .Q(n83) );
  INV3 U544 ( .A(n191), .Q(n287) );
  INV3 U545 ( .A(n141), .Q(n281) );
  INV3 U546 ( .A(n209), .Q(n289) );
  NAND22 U547 ( .A(n291), .B(n224), .Q(n26) );
  INV0 U548 ( .A(n223), .Q(n291) );
  INV3 U549 ( .A(n124), .Q(n122) );
  INV3 U550 ( .A(n192), .Q(n190) );
  AOI210 U551 ( .A(n147), .B(n281), .C(n140), .Q(n138) );
  INV3 U552 ( .A(n142), .Q(n140) );
  INV3 U553 ( .A(n86), .Q(n84) );
  XNR21 U554 ( .A(n6), .B(n49), .Q(SUM[29]) );
  NAND22 U555 ( .A(n288), .B(n203), .Q(n23) );
  INV3 U556 ( .A(n202), .Q(n288) );
  NAND22 U557 ( .A(n276), .B(n97), .Q(n11) );
  NAND22 U558 ( .A(n279), .B(n124), .Q(n14) );
  NAND22 U559 ( .A(n274), .B(n79), .Q(n9) );
  INV3 U560 ( .A(n78), .Q(n274) );
  INV0 U561 ( .A(n152), .Q(n282) );
  NAND22 U562 ( .A(n286), .B(n185), .Q(n21) );
  INV3 U563 ( .A(n184), .Q(n286) );
  NAND22 U564 ( .A(n277), .B(n106), .Q(n12) );
  NAND22 U565 ( .A(n281), .B(n142), .Q(n16) );
  INV0 U566 ( .A(n147), .Q(n145) );
  NAND22 U567 ( .A(n278), .B(n117), .Q(n13) );
  INV0 U568 ( .A(n116), .Q(n278) );
  NAND22 U569 ( .A(n272), .B(n59), .Q(n7) );
  INV3 U570 ( .A(n58), .Q(n272) );
  NAND22 U571 ( .A(n285), .B(n174), .Q(n20) );
  INV0 U572 ( .A(n171), .Q(n285) );
  NAND20 U573 ( .A(n289), .B(n210), .Q(n24) );
  NAND21 U574 ( .A(n296), .B(n259), .Q(n31) );
  NAND22 U575 ( .A(n295), .B(n253), .Q(n30) );
  NAND22 U576 ( .A(n292), .B(n232), .Q(n27) );
  INV0 U577 ( .A(n231), .Q(n292) );
  INV3 U578 ( .A(n253), .Q(n251) );
  XOR20 U579 ( .A(n268), .B(n33), .Q(SUM[2]) );
  NOR21 U580 ( .A(B[29]), .B(A[29]), .Q(n47) );
  NOR22 U581 ( .A(B[20]), .B(A[20]), .Q(n134) );
  XOR21 U582 ( .A(n4), .B(n37), .Q(SUM[31]) );
  NAND22 U583 ( .A(n269), .B(n36), .Q(n4) );
  NAND22 U584 ( .A(A[31]), .B(B[31]), .Q(n36) );
  NAND20 U585 ( .A(n299), .B(n268), .Q(n34) );
  INV2 U586 ( .A(n267), .Q(n299) );
  INV3 U587 ( .A(n40), .Q(n38) );
  INV3 U588 ( .A(n35), .Q(n269) );
  NOR21 U589 ( .A(B[31]), .B(A[31]), .Q(n35) );
  BUF2 U590 ( .A(A[0]), .Q(SUM[0]) );
  LOGIC0 U591 ( .Q(n39) );
  OAI211 U592 ( .A(n70), .B(n425), .C(n71), .Q(n69) );
  NAND22 U593 ( .A(A[7]), .B(B[7]), .Q(n239) );
  NOR23 U594 ( .A(B[3]), .B(A[3]), .Q(n261) );
  OAI211 U595 ( .A(n43), .B(n415), .C(n44), .Q(n42) );
  CLKIN0 U596 ( .A(n164), .Q(n284) );
  NOR22 U597 ( .A(B[5]), .B(A[5]), .Q(n252) );
  NOR22 U598 ( .A(n160), .B(n194), .Q(n158) );
  NAND24 U599 ( .A(n178), .B(n162), .Q(n160) );
  AOI212 U600 ( .A(n226), .B(n158), .C(n159), .Q(n1) );
  AOI210 U601 ( .A(n2), .B(n52), .C(n53), .Q(n51) );
  AOI210 U602 ( .A(n2), .B(n45), .C(n46), .Q(n44) );
  AOI211 U603 ( .A(n2), .B(n72), .C(n73), .Q(n71) );
  NOR23 U604 ( .A(B[8]), .B(A[8]), .Q(n231) );
  NOR20 U605 ( .A(B[1]), .B(A[1]), .Q(n267) );
endmodule


module sqroot_seq_NBITS32_DW01_sub_7 ( A, B, CI, DIFF, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n68, n69, n70, n71, n72, n73, n74, n75,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n106, n107,
         n108, n109, n110, n111, n112, n113, n116, n117, n118, n119, n120,
         n122, n123, n124, n125, n126, n127, n128, n129, n132, n133, n134,
         n135, n136, n137, n138, n140, n141, n142, n143, n144, n145, n146,
         n147, n152, n153, n154, n155, n156, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n174, n175,
         n176, n177, n178, n179, n180, n181, n184, n185, n186, n187, n188,
         n190, n191, n192, n193, n194, n195, n196, n197, n200, n201, n202,
         n203, n204, n205, n206, n208, n209, n210, n211, n212, n213, n214,
         n215, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n239, n240, n241, n242,
         n243, n244, n247, n248, n249, n251, n252, n253, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502;

  XNR22 U11 ( .A(n5), .B(n42), .Q(DIFF[29]) );
  XNR22 U19 ( .A(n6), .B(n49), .Q(DIFF[28]) );
  OAI212 U20 ( .A(n43), .B(n502), .C(n44), .Q(n42) );
  NOR24 U23 ( .A(n47), .B(n54), .Q(n45) );
  OAI212 U24 ( .A(n47), .B(n55), .C(n48), .Q(n46) );
  AOI212 U36 ( .A(n73), .B(n56), .C(n57), .Q(n55) );
  OAI212 U38 ( .A(n68), .B(n58), .C(n59), .Q(n57) );
  OAI212 U44 ( .A(n61), .B(n453), .C(n62), .Q(n60) );
  OAI212 U56 ( .A(n70), .B(n453), .C(n71), .Q(n69) );
  OAI212 U64 ( .A(n86), .B(n78), .C(n79), .Q(n73) );
  OAI212 U70 ( .A(n81), .B(n502), .C(n82), .Q(n80) );
  AOI212 U72 ( .A(n488), .B(n83), .C(n84), .Q(n82) );
  OAI212 U80 ( .A(n88), .B(n452), .C(n89), .Q(n87) );
  OAI212 U84 ( .A(n92), .B(n127), .C(n93), .Q(n2) );
  OAI212 U88 ( .A(n106), .B(n96), .C(n97), .Q(n95) );
  OAI212 U94 ( .A(n99), .B(n502), .C(n100), .Q(n98) );
  OAI212 U98 ( .A(n103), .B(n113), .C(n106), .Q(n102) );
  OAI212 U106 ( .A(n108), .B(n502), .C(n109), .Q(n107) );
  OAI212 U114 ( .A(n124), .B(n116), .C(n117), .Q(n111) );
  OAI212 U120 ( .A(n119), .B(n502), .C(n120), .Q(n118) );
  AOI212 U136 ( .A(n147), .B(n132), .C(n133), .Q(n127) );
  OAI212 U138 ( .A(n142), .B(n134), .C(n135), .Q(n133) );
  OAI212 U144 ( .A(n137), .B(n502), .C(n138), .Q(n136) );
  OAI212 U154 ( .A(n144), .B(n502), .C(n145), .Q(n143) );
  OAI212 U162 ( .A(n156), .B(n152), .C(n153), .Q(n147) );
  OAI212 U168 ( .A(n155), .B(n502), .C(n156), .Q(n154) );
  AOI212 U174 ( .A(n226), .B(n158), .C(n159), .Q(n1) );
  OAI212 U176 ( .A(n160), .B(n195), .C(n161), .Q(n159) );
  AOI212 U178 ( .A(n179), .B(n162), .C(n163), .Q(n161) );
  NOR24 U179 ( .A(n164), .B(n171), .Q(n162) );
  OAI212 U180 ( .A(n174), .B(n164), .C(n165), .Q(n163) );
  NOR24 U183 ( .A(A[15]), .B(n313), .Q(n164) );
  OAI212 U190 ( .A(n171), .B(n181), .C(n174), .Q(n170) );
  NOR24 U195 ( .A(A[14]), .B(n314), .Q(n171) );
  XNR22 U197 ( .A(n21), .B(n186), .Q(DIFF[13]) );
  NOR24 U205 ( .A(n184), .B(n191), .Q(n178) );
  OAI212 U206 ( .A(n192), .B(n184), .C(n185), .Q(n179) );
  NOR24 U209 ( .A(A[13]), .B(n315), .Q(n184) );
  OAI212 U212 ( .A(n187), .B(n481), .C(n188), .Q(n186) );
  AOI212 U228 ( .A(n215), .B(n200), .C(n201), .Q(n195) );
  OAI212 U230 ( .A(n210), .B(n202), .C(n203), .Q(n201) );
  NOR24 U233 ( .A(A[11]), .B(n317), .Q(n202) );
  XNR22 U235 ( .A(n24), .B(n211), .Q(DIFF[10]) );
  OAI212 U236 ( .A(n205), .B(n498), .C(n206), .Q(n204) );
  OAI212 U246 ( .A(n212), .B(n481), .C(n213), .Q(n211) );
  OAI212 U254 ( .A(n224), .B(n220), .C(n221), .Q(n215) );
  OAI212 U260 ( .A(n223), .B(n498), .C(n224), .Q(n222) );
  AOI212 U269 ( .A(n242), .B(n229), .C(n230), .Q(n228) );
  OAI212 U271 ( .A(n239), .B(n231), .C(n232), .Q(n230) );
  NOR24 U274 ( .A(A[7]), .B(n321), .Q(n231) );
  AOI212 U277 ( .A(n435), .B(n234), .C(n235), .Q(n233) );
  OAI212 U279 ( .A(n244), .B(n236), .C(n239), .Q(n235) );
  NOR24 U284 ( .A(A[6]), .B(n322), .Q(n236) );
  XOR22 U286 ( .A(n29), .B(n249), .Q(DIFF[5]) );
  OAI212 U293 ( .A(n253), .B(n247), .C(n248), .Q(n242) );
  XNR22 U298 ( .A(n30), .B(n435), .Q(DIFF[4]) );
  XNR22 U306 ( .A(n31), .B(n260), .Q(DIFF[3]) );
  AOI212 U308 ( .A(n264), .B(n256), .C(n257), .Q(n255) );
  OAI212 U310 ( .A(n262), .B(n258), .C(n259), .Q(n257) );
  NOR24 U313 ( .A(A[3]), .B(n325), .Q(n258) );
  OAI212 U323 ( .A(n267), .B(n265), .C(n266), .Q(n264) );
  CLKIN6 U364 ( .A(n41), .Q(n5) );
  AOI211 U365 ( .A(n42), .B(n38), .C(n39), .Q(n37) );
  CLKIN6 U366 ( .A(A[29]), .Q(n41) );
  NAND24 U367 ( .A(n433), .B(n434), .Q(DIFF[20]) );
  INV6 U368 ( .A(n125), .Q(n431) );
  CLKIN8 U369 ( .A(B[5]), .Q(n323) );
  NAND26 U370 ( .A(n501), .B(n228), .Q(n226) );
  OAI211 U371 ( .A(n253), .B(n247), .C(n248), .Q(n451) );
  NAND23 U372 ( .A(n324), .B(A[4]), .Q(n253) );
  CLKIN3 U373 ( .A(n154), .Q(n482) );
  NOR23 U374 ( .A(A[5]), .B(n323), .Q(n247) );
  NOR24 U375 ( .A(A[5]), .B(n323), .Q(n486) );
  NOR24 U376 ( .A(A[1]), .B(n327), .Q(n265) );
  CLKIN4 U377 ( .A(B[1]), .Q(n327) );
  CLKIN3 U378 ( .A(n136), .Q(n477) );
  NAND23 U379 ( .A(n154), .B(n17), .Q(n484) );
  NOR22 U380 ( .A(A[26]), .B(n302), .Q(n65) );
  XNR22 U381 ( .A(n9), .B(n80), .Q(DIFF[25]) );
  CLKIN8 U382 ( .A(n502), .Q(n492) );
  NOR23 U383 ( .A(A[9]), .B(n319), .Q(n220) );
  NAND26 U384 ( .A(n471), .B(n168), .Q(n166) );
  AOI211 U385 ( .A(n197), .B(n169), .C(n170), .Q(n168) );
  AOI211 U386 ( .A(n111), .B(n94), .C(n95), .Q(n93) );
  NAND23 U387 ( .A(n318), .B(A[10]), .Q(n210) );
  NAND22 U388 ( .A(n312), .B(A[16]), .Q(n156) );
  NAND24 U389 ( .A(n492), .B(n128), .Q(n493) );
  INV3 U390 ( .A(B[4]), .Q(n324) );
  NAND22 U391 ( .A(n443), .B(n444), .Q(DIFF[12]) );
  NAND22 U392 ( .A(n441), .B(n442), .Q(n444) );
  NAND22 U393 ( .A(n481), .B(n494), .Q(n497) );
  INV12 U394 ( .A(n498), .Q(n470) );
  CLKIN4 U395 ( .A(n225), .Q(n495) );
  NAND23 U396 ( .A(n326), .B(A[2]), .Q(n262) );
  NAND22 U397 ( .A(n125), .B(n14), .Q(n433) );
  NAND23 U398 ( .A(n431), .B(n432), .Q(n434) );
  INV3 U399 ( .A(n14), .Q(n432) );
  NAND23 U400 ( .A(n493), .B(n127), .Q(n125) );
  NAND26 U401 ( .A(n484), .B(n485), .Q(DIFF[17]) );
  INV3 U402 ( .A(n492), .Q(n452) );
  INV3 U403 ( .A(n178), .Q(n180) );
  CLKIN10 U404 ( .A(n166), .Q(n473) );
  NAND23 U405 ( .A(n19), .B(n166), .Q(n474) );
  CLKBU12 U406 ( .A(n500), .Q(n435) );
  INV6 U407 ( .A(n255), .Q(n500) );
  INV2 U408 ( .A(n296), .Q(n436) );
  INV3 U409 ( .A(n261), .Q(n296) );
  NOR23 U410 ( .A(A[2]), .B(n326), .Q(n261) );
  NOR22 U411 ( .A(n65), .B(n74), .Q(n63) );
  NAND21 U412 ( .A(n302), .B(A[26]), .Q(n68) );
  NAND24 U413 ( .A(n316), .B(A[12]), .Q(n192) );
  NAND26 U414 ( .A(n479), .B(n480), .Q(DIFF[19]) );
  NAND22 U415 ( .A(n16), .B(n143), .Q(n439) );
  NAND24 U416 ( .A(n437), .B(n438), .Q(n440) );
  NAND24 U417 ( .A(n439), .B(n440), .Q(DIFF[18]) );
  INV1 U418 ( .A(n16), .Q(n437) );
  INV3 U419 ( .A(n143), .Q(n438) );
  CLKIN3 U420 ( .A(n141), .Q(n280) );
  NOR23 U421 ( .A(n134), .B(n141), .Q(n132) );
  NAND23 U422 ( .A(n136), .B(n15), .Q(n479) );
  NAND24 U423 ( .A(n469), .B(n470), .Q(n471) );
  NAND21 U424 ( .A(n296), .B(n262), .Q(n32) );
  INV3 U425 ( .A(n209), .Q(n288) );
  NOR22 U426 ( .A(n258), .B(n261), .Q(n256) );
  CLKIN3 U427 ( .A(n146), .Q(n144) );
  NOR22 U428 ( .A(n152), .B(n155), .Q(n146) );
  INV2 U429 ( .A(n127), .Q(n129) );
  INV3 U430 ( .A(B[22]), .Q(n306) );
  NOR22 U431 ( .A(A[4]), .B(n324), .Q(n252) );
  INV3 U432 ( .A(n27), .Q(n476) );
  INV3 U433 ( .A(B[15]), .Q(n313) );
  INV3 U434 ( .A(B[12]), .Q(n316) );
  NOR23 U435 ( .A(A[12]), .B(n316), .Q(n191) );
  INV3 U436 ( .A(n167), .Q(n469) );
  INV3 U437 ( .A(B[17]), .Q(n311) );
  NOR21 U438 ( .A(A[18]), .B(n310), .Q(n141) );
  INV3 U439 ( .A(B[19]), .Q(n309) );
  INV3 U440 ( .A(B[18]), .Q(n310) );
  INV3 U441 ( .A(B[21]), .Q(n307) );
  INV3 U442 ( .A(n227), .Q(n499) );
  NOR21 U443 ( .A(n78), .B(n85), .Q(n72) );
  NOR21 U444 ( .A(A[24]), .B(n304), .Q(n85) );
  NOR23 U445 ( .A(A[10]), .B(n318), .Q(n209) );
  INV3 U446 ( .A(B[16]), .Q(n312) );
  NOR23 U447 ( .A(A[17]), .B(n311), .Q(n152) );
  NOR22 U448 ( .A(A[19]), .B(n309), .Q(n134) );
  NOR21 U449 ( .A(n103), .B(n112), .Q(n101) );
  NAND23 U450 ( .A(n214), .B(n200), .Q(n194) );
  NOR21 U451 ( .A(A[27]), .B(n301), .Q(n58) );
  NOR22 U452 ( .A(n92), .B(n126), .Q(n3) );
  AOI211 U453 ( .A(n488), .B(n52), .C(n53), .Q(n51) );
  INV3 U454 ( .A(n204), .Q(n448) );
  CLKIN3 U455 ( .A(n175), .Q(n455) );
  NOR22 U456 ( .A(A[16]), .B(n312), .Q(n155) );
  INV3 U457 ( .A(n118), .Q(n460) );
  NOR22 U458 ( .A(A[22]), .B(n306), .Q(n103) );
  INV3 U459 ( .A(n223), .Q(n290) );
  XOR21 U460 ( .A(n4), .B(n37), .Q(DIFF[30]) );
  INV3 U461 ( .A(n28), .Q(n458) );
  NAND24 U462 ( .A(n467), .B(n468), .Q(DIFF[9]) );
  NAND24 U463 ( .A(n465), .B(n466), .Q(n468) );
  NAND22 U464 ( .A(n22), .B(n193), .Q(n443) );
  INV2 U465 ( .A(n22), .Q(n441) );
  INV4 U466 ( .A(n193), .Q(n442) );
  CLKIN6 U467 ( .A(B[9]), .Q(n319) );
  NAND21 U468 ( .A(n294), .B(n253), .Q(n30) );
  INV2 U469 ( .A(n213), .Q(n445) );
  INV2 U470 ( .A(n215), .Q(n213) );
  BUF2 U471 ( .A(n202), .Q(n446) );
  NAND22 U472 ( .A(n23), .B(n204), .Q(n449) );
  NAND24 U473 ( .A(n447), .B(n448), .Q(n450) );
  NAND24 U474 ( .A(n449), .B(n450), .Q(DIFF[11]) );
  INV3 U475 ( .A(n23), .Q(n447) );
  INV3 U476 ( .A(n451), .Q(n244) );
  INV4 U477 ( .A(n492), .Q(n453) );
  NAND22 U478 ( .A(n20), .B(n175), .Q(n456) );
  NAND24 U479 ( .A(n454), .B(n455), .Q(n457) );
  NAND28 U480 ( .A(n456), .B(n457), .Q(DIFF[14]) );
  INV3 U481 ( .A(n20), .Q(n454) );
  NAND22 U482 ( .A(n284), .B(n174), .Q(n20) );
  OAI211 U483 ( .A(n50), .B(n502), .C(n51), .Q(n49) );
  INV1 U484 ( .A(n197), .Q(n489) );
  XOR21 U485 ( .A(n32), .B(n263), .Q(DIFF[2]) );
  XNR22 U486 ( .A(n458), .B(n240), .Q(DIFF[6]) );
  NAND28 U487 ( .A(n472), .B(n473), .Q(n475) );
  NOR24 U488 ( .A(n231), .B(n236), .Q(n229) );
  NAND22 U489 ( .A(n222), .B(n25), .Q(n467) );
  NAND24 U490 ( .A(n496), .B(n497), .Q(DIFF[8]) );
  NAND22 U491 ( .A(n295), .B(n259), .Q(n31) );
  NAND21 U492 ( .A(n26), .B(n495), .Q(n496) );
  INV3 U493 ( .A(B[25]), .Q(n303) );
  NAND21 U494 ( .A(n303), .B(A[25]), .Q(n79) );
  NAND22 U495 ( .A(n13), .B(n118), .Q(n461) );
  NAND24 U496 ( .A(n459), .B(n460), .Q(n462) );
  NAND24 U497 ( .A(n461), .B(n462), .Q(DIFF[21]) );
  INV3 U498 ( .A(n13), .Q(n459) );
  XNR22 U499 ( .A(n10), .B(n87), .Q(DIFF[24]) );
  OAI211 U500 ( .A(n35), .B(n37), .C(n36), .Q(n34) );
  NOR22 U501 ( .A(A[9]), .B(n319), .Q(n463) );
  OAI211 U502 ( .A(n267), .B(n265), .C(n266), .Q(n464) );
  NAND28 U503 ( .A(n474), .B(n475), .Q(DIFF[15]) );
  NAND24 U504 ( .A(n196), .B(n470), .Q(n491) );
  INV3 U505 ( .A(n222), .Q(n465) );
  INV2 U506 ( .A(n25), .Q(n466) );
  NAND21 U507 ( .A(n289), .B(n221), .Q(n25) );
  CLKIN6 U508 ( .A(n19), .Q(n472) );
  NAND26 U509 ( .A(n491), .B(n489), .Q(n193) );
  XNR22 U510 ( .A(n476), .B(n233), .Q(DIFF[7]) );
  NAND26 U511 ( .A(n477), .B(n478), .Q(n480) );
  CLKIN6 U512 ( .A(n15), .Q(n478) );
  INV2 U513 ( .A(n241), .Q(n243) );
  NAND26 U514 ( .A(n320), .B(A[8]), .Q(n224) );
  INV3 U515 ( .A(n54), .Q(n52) );
  CLKIN3 U516 ( .A(n55), .Q(n53) );
  INV6 U517 ( .A(n495), .Q(n481) );
  INV4 U518 ( .A(n226), .Q(n225) );
  NAND24 U519 ( .A(n241), .B(n229), .Q(n227) );
  CLKBU15 U520 ( .A(n1), .Q(n502) );
  NAND21 U521 ( .A(n282), .B(n156), .Q(n18) );
  XOR21 U522 ( .A(n267), .B(n33), .Q(DIFF[1]) );
  XNR22 U523 ( .A(n7), .B(n60), .Q(DIFF[27]) );
  NOR24 U524 ( .A(n486), .B(n252), .Q(n241) );
  NAND21 U525 ( .A(n3), .B(n83), .Q(n81) );
  NAND21 U526 ( .A(n285), .B(n185), .Q(n21) );
  AOI210 U527 ( .A(n197), .B(n178), .C(n179), .Q(n177) );
  OAI212 U528 ( .A(n436), .B(n263), .C(n262), .Q(n260) );
  NAND26 U529 ( .A(n482), .B(n483), .Q(n485) );
  CLKIN6 U530 ( .A(n17), .Q(n483) );
  NAND24 U531 ( .A(n500), .B(n499), .Q(n501) );
  BUF2 U532 ( .A(n258), .Q(n487) );
  BUF12 U533 ( .A(n2), .Q(n488) );
  INV1 U534 ( .A(n265), .Q(n297) );
  XNR22 U535 ( .A(n11), .B(n98), .Q(DIFF[23]) );
  NAND22 U536 ( .A(n196), .B(n169), .Q(n167) );
  NOR21 U537 ( .A(n171), .B(n180), .Q(n169) );
  NOR22 U538 ( .A(A[25]), .B(n303), .Q(n78) );
  INV2 U539 ( .A(n179), .Q(n181) );
  NAND22 U540 ( .A(n325), .B(A[3]), .Q(n259) );
  INV2 U541 ( .A(n464), .Q(n263) );
  OAI211 U542 ( .A(n65), .B(n75), .C(n68), .Q(n64) );
  NOR23 U543 ( .A(n58), .B(n65), .Q(n56) );
  INV1 U544 ( .A(n65), .Q(n272) );
  XNR22 U545 ( .A(n8), .B(n69), .Q(DIFF[26]) );
  XNR22 U546 ( .A(n12), .B(n107), .Q(DIFF[22]) );
  CLKIN1 U547 ( .A(B[24]), .Q(n304) );
  NAND22 U548 ( .A(n313), .B(A[15]), .Q(n165) );
  AOI212 U549 ( .A(n435), .B(n294), .C(n251), .Q(n249) );
  NAND20 U550 ( .A(n305), .B(A[23]), .Q(n490) );
  NAND22 U551 ( .A(n305), .B(A[23]), .Q(n97) );
  INV2 U552 ( .A(B[23]), .Q(n305) );
  CLKIN6 U553 ( .A(B[3]), .Q(n325) );
  CLKIN6 U554 ( .A(B[2]), .Q(n326) );
  CLKBU15 U555 ( .A(n225), .Q(n498) );
  NAND22 U556 ( .A(n128), .B(n101), .Q(n99) );
  INV1 U557 ( .A(n110), .Q(n112) );
  NAND21 U558 ( .A(n307), .B(A[21]), .Q(n117) );
  XOR21 U559 ( .A(n18), .B(n502), .Q(DIFF[16]) );
  NAND22 U560 ( .A(n146), .B(n132), .Q(n126) );
  NAND20 U561 ( .A(n290), .B(n224), .Q(n26) );
  INV2 U562 ( .A(n26), .Q(n494) );
  NAND21 U563 ( .A(n128), .B(n110), .Q(n108) );
  NOR22 U564 ( .A(n116), .B(n123), .Q(n110) );
  CLKIN1 U565 ( .A(n123), .Q(n278) );
  CLKIN6 U566 ( .A(B[0]), .Q(n328) );
  NAND24 U567 ( .A(n327), .B(A[1]), .Q(n266) );
  CLKIN3 U568 ( .A(n126), .Q(n128) );
  NAND20 U569 ( .A(n196), .B(n286), .Q(n187) );
  INV0 U570 ( .A(n191), .Q(n286) );
  INV0 U571 ( .A(n253), .Q(n251) );
  INV6 U572 ( .A(B[6]), .Q(n322) );
  OAI212 U573 ( .A(n176), .B(n498), .C(n177), .Q(n175) );
  XNR20 U574 ( .A(n328), .B(A[0]), .Q(DIFF[0]) );
  NAND20 U575 ( .A(n146), .B(n280), .Q(n137) );
  NAND20 U576 ( .A(n214), .B(n288), .Q(n205) );
  NOR24 U577 ( .A(A[0]), .B(n328), .Q(n267) );
  NOR22 U578 ( .A(n160), .B(n194), .Q(n158) );
  NAND20 U579 ( .A(n3), .B(n72), .Q(n70) );
  AOI210 U580 ( .A(n488), .B(n72), .C(n73), .Q(n71) );
  INV0 U581 ( .A(n171), .Q(n284) );
  NAND20 U582 ( .A(n280), .B(n142), .Q(n16) );
  AOI211 U583 ( .A(n488), .B(n63), .C(n64), .Q(n62) );
  CLKIN2 U584 ( .A(n73), .Q(n75) );
  NAND21 U585 ( .A(n3), .B(n45), .Q(n43) );
  AOI211 U586 ( .A(n488), .B(n45), .C(n46), .Q(n44) );
  NOR23 U587 ( .A(n202), .B(n209), .Q(n200) );
  NAND21 U588 ( .A(n270), .B(n48), .Q(n6) );
  NAND20 U589 ( .A(n272), .B(n68), .Q(n8) );
  INV1 U590 ( .A(n3), .Q(n88) );
  NAND20 U591 ( .A(n83), .B(n86), .Q(n10) );
  NAND23 U592 ( .A(n322), .B(A[6]), .Q(n239) );
  CLKIN3 U593 ( .A(B[27]), .Q(n301) );
  INV1 U594 ( .A(n488), .Q(n89) );
  NOR22 U595 ( .A(n96), .B(n103), .Q(n94) );
  CLKIN0 U596 ( .A(n116), .Q(n277) );
  CLKIN0 U597 ( .A(n103), .Q(n276) );
  CLKIN0 U598 ( .A(n210), .Q(n208) );
  CLKIN0 U599 ( .A(n142), .Q(n140) );
  CLKIN0 U600 ( .A(n236), .Q(n292) );
  NAND20 U601 ( .A(n286), .B(n192), .Q(n22) );
  INV2 U602 ( .A(n72), .Q(n74) );
  CLKIN0 U603 ( .A(n164), .Q(n283) );
  INV0 U604 ( .A(n47), .Q(n270) );
  INV0 U605 ( .A(n487), .Q(n295) );
  NOR22 U606 ( .A(A[23]), .B(n305), .Q(n96) );
  NAND21 U607 ( .A(n315), .B(A[13]), .Q(n185) );
  NAND21 U608 ( .A(n304), .B(A[24]), .Q(n86) );
  NAND21 U609 ( .A(n308), .B(A[20]), .Q(n124) );
  NAND21 U610 ( .A(n306), .B(A[22]), .Q(n106) );
  NAND20 U611 ( .A(n300), .B(A[28]), .Q(n48) );
  NAND20 U612 ( .A(n301), .B(A[27]), .Q(n59) );
  CLKIN3 U613 ( .A(B[28]), .Q(n300) );
  NOR24 U614 ( .A(A[8]), .B(n320), .Q(n223) );
  NAND22 U615 ( .A(n3), .B(n52), .Q(n50) );
  INV3 U616 ( .A(n194), .Q(n196) );
  AOI210 U617 ( .A(n129), .B(n110), .C(n111), .Q(n109) );
  NAND22 U618 ( .A(n72), .B(n56), .Q(n54) );
  NAND22 U619 ( .A(n178), .B(n162), .Q(n160) );
  NAND22 U620 ( .A(n110), .B(n94), .Q(n92) );
  NAND22 U621 ( .A(n3), .B(n63), .Q(n61) );
  NAND20 U622 ( .A(n196), .B(n178), .Q(n176) );
  NAND22 U623 ( .A(n128), .B(n278), .Q(n119) );
  NAND22 U624 ( .A(n297), .B(n266), .Q(n33) );
  NAND22 U625 ( .A(n292), .B(n239), .Q(n28) );
  NAND22 U626 ( .A(n268), .B(n36), .Q(n4) );
  INV3 U627 ( .A(n35), .Q(n268) );
  INV3 U628 ( .A(n155), .Q(n282) );
  NAND22 U629 ( .A(n283), .B(n165), .Q(n19) );
  NAND22 U630 ( .A(n273), .B(n79), .Q(n9) );
  INV3 U631 ( .A(n78), .Q(n273) );
  NAND22 U632 ( .A(n277), .B(n117), .Q(n13) );
  NOR22 U633 ( .A(n463), .B(n223), .Q(n214) );
  INV0 U634 ( .A(n463), .Q(n289) );
  NAND22 U635 ( .A(n278), .B(n124), .Q(n14) );
  NAND22 U636 ( .A(n279), .B(n135), .Q(n15) );
  INV0 U637 ( .A(n134), .Q(n279) );
  INV0 U638 ( .A(n184), .Q(n285) );
  NAND22 U639 ( .A(n287), .B(n203), .Q(n23) );
  INV0 U640 ( .A(n446), .Q(n287) );
  NAND22 U641 ( .A(n288), .B(n210), .Q(n24) );
  INV0 U642 ( .A(n214), .Q(n212) );
  INV0 U643 ( .A(n147), .Q(n145) );
  NAND22 U644 ( .A(n275), .B(n490), .Q(n11) );
  INV3 U645 ( .A(n96), .Q(n275) );
  NAND22 U646 ( .A(n271), .B(n59), .Q(n7) );
  INV3 U647 ( .A(n58), .Q(n271) );
  NAND22 U648 ( .A(n276), .B(n106), .Q(n12) );
  NAND22 U649 ( .A(n281), .B(n153), .Q(n17) );
  INV0 U650 ( .A(n152), .Q(n281) );
  NAND22 U651 ( .A(n291), .B(n232), .Q(n27) );
  INV0 U652 ( .A(n231), .Q(n291) );
  NAND20 U653 ( .A(n293), .B(n248), .Q(n29) );
  INV3 U654 ( .A(n85), .Q(n83) );
  INV3 U655 ( .A(n86), .Q(n84) );
  AOI211 U656 ( .A(n129), .B(n101), .C(n102), .Q(n100) );
  INV0 U657 ( .A(n111), .Q(n113) );
  AOI210 U658 ( .A(n197), .B(n286), .C(n190), .Q(n188) );
  INV3 U659 ( .A(n192), .Q(n190) );
  AOI211 U660 ( .A(n129), .B(n278), .C(n122), .Q(n120) );
  INV3 U661 ( .A(n124), .Q(n122) );
  AOI210 U662 ( .A(n147), .B(n280), .C(n140), .Q(n138) );
  NOR20 U663 ( .A(n236), .B(n243), .Q(n234) );
  INV3 U664 ( .A(n252), .Q(n294) );
  XNR21 U665 ( .A(A[31]), .B(n34), .Q(DIFF[31]) );
  NOR21 U666 ( .A(A[28]), .B(n300), .Q(n47) );
  INV3 U667 ( .A(n41), .Q(n39) );
  NOR23 U668 ( .A(A[21]), .B(n307), .Q(n116) );
  NOR21 U669 ( .A(A[20]), .B(n308), .Q(n123) );
  NAND22 U670 ( .A(n310), .B(A[18]), .Q(n142) );
  NAND22 U671 ( .A(n314), .B(A[14]), .Q(n174) );
  NAND22 U672 ( .A(n317), .B(A[11]), .Q(n203) );
  NAND22 U673 ( .A(n321), .B(A[7]), .Q(n232) );
  NAND22 U674 ( .A(n311), .B(A[17]), .Q(n153) );
  NAND22 U675 ( .A(n309), .B(A[19]), .Q(n135) );
  NAND22 U676 ( .A(n319), .B(A[9]), .Q(n221) );
  CLKIN3 U677 ( .A(B[20]), .Q(n308) );
  INV3 U678 ( .A(B[26]), .Q(n302) );
  NOR21 U679 ( .A(A[30]), .B(n298), .Q(n35) );
  NAND22 U680 ( .A(n298), .B(A[30]), .Q(n36) );
  INV3 U681 ( .A(B[30]), .Q(n298) );
  LOGIC1 U682 ( .Q(n38) );
  AOI211 U683 ( .A(n435), .B(n241), .C(n242), .Q(n240) );
  NAND22 U684 ( .A(n323), .B(A[5]), .Q(n248) );
  INV3 U685 ( .A(n486), .Q(n293) );
  AOI210 U686 ( .A(n445), .B(n288), .C(n208), .Q(n206) );
  CLKIN2 U687 ( .A(n195), .Q(n197) );
  CLKIN6 U688 ( .A(B[7]), .Q(n321) );
  CLKIN6 U689 ( .A(B[8]), .Q(n320) );
  CLKIN6 U690 ( .A(B[10]), .Q(n318) );
  CLKIN6 U691 ( .A(B[11]), .Q(n317) );
  CLKIN6 U692 ( .A(B[13]), .Q(n315) );
  CLKIN6 U693 ( .A(B[14]), .Q(n314) );
endmodule


module sqroot_seq_NBITS32 ( arg, roundup, clk, nRst, start, sqroot, ready );
  input [31:0] arg;
  output [16:0] sqroot;
  input roundup, clk, nRst, start;
  output ready;
  wire   n_Logic0_, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, N40, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51,
         N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65,
         N66, N67, N68, N69, N70, N71, N72, N73, N74, n37, n38, n39, n42, n4,
         n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65, n66, n212, n213, N99, N98,
         N97, N96, N95, N94, N93, N92, N91, N90, N89, N120, N119, N118, N117,
         N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, N106,
         N105, N104, N103, N102, N101, N100, n215, n216, n217, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n232,
         n233, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n249, n250, n251, n252, n253, n254, n256, n258,
         n260, n261, n262, n264, n265, n266, n267, n268, n269, n270, n273,
         n274, n275, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472;
  wire   [2:0] state_reg;
  wire   [31:17] root_reg;
  wire   [30:0] delta_reg;
  wire   [31:0] res_reg;
  wire   [31:0] root_next;
  wire   [30:6] delta_next;
  wire   [30:0] res_next;
  wire   [31:0] fuo_if_res;
  wire   [31:0] fuo_if_root;
  wire   [31:0] fuo_round;

  DFC3 delta_reg_reg_10_ ( .D(delta_next[10]), .C(clk), .RN(nRst), .Q(
        delta_reg[10]), .QN(n62) );
  DFC3 delta_reg_reg_30_ ( .D(delta_next[30]), .C(clk), .RN(nRst), .Q(
        delta_reg[30]), .QN(n42) );
  DFC3 delta_reg_reg_28_ ( .D(delta_next[28]), .C(clk), .RN(nRst), .Q(
        delta_reg[28]), .QN(n44) );
  DFC3 delta_reg_reg_26_ ( .D(delta_next[26]), .C(clk), .RN(nRst), .Q(
        delta_reg[26]), .QN(n46) );
  DFC3 delta_reg_reg_24_ ( .D(delta_next[24]), .C(clk), .RN(nRst), .Q(
        delta_reg[24]), .QN(n48) );
  DFC3 delta_reg_reg_22_ ( .D(delta_next[22]), .C(clk), .RN(nRst), .Q(
        delta_reg[22]), .QN(n50) );
  DFC3 delta_reg_reg_20_ ( .D(delta_next[20]), .C(clk), .RN(nRst), .Q(
        delta_reg[20]), .QN(n52) );
  DFC3 delta_reg_reg_18_ ( .D(delta_next[18]), .C(clk), .RN(nRst), .Q(
        delta_reg[18]), .QN(n54) );
  DFC3 delta_reg_reg_16_ ( .D(delta_next[16]), .C(clk), .RN(nRst), .Q(
        delta_reg[16]), .QN(n56) );
  DFC3 delta_reg_reg_14_ ( .D(delta_next[14]), .C(clk), .RN(nRst), .Q(
        delta_reg[14]), .QN(n58) );
  DFC3 delta_reg_reg_12_ ( .D(delta_next[12]), .C(clk), .RN(nRst), .Q(
        delta_reg[12]), .QN(n60) );
  DFC3 delta_reg_reg_8_ ( .D(delta_next[8]), .C(clk), .RN(nRst), .Q(
        delta_reg[8]), .QN(n64) );
  DFC3 delta_reg_reg_27_ ( .D(delta_next[27]), .C(clk), .RN(nRst), .Q(
        delta_reg[27]), .QN(n45) );
  DFC3 delta_reg_reg_25_ ( .D(delta_next[25]), .C(clk), .RN(nRst), .Q(
        delta_reg[25]), .QN(n47) );
  DFC3 delta_reg_reg_23_ ( .D(delta_next[23]), .C(clk), .RN(nRst), .Q(
        delta_reg[23]), .QN(n49) );
  DFC3 delta_reg_reg_21_ ( .D(delta_next[21]), .C(clk), .RN(nRst), .Q(
        delta_reg[21]), .QN(n51) );
  DFC3 delta_reg_reg_19_ ( .D(delta_next[19]), .C(clk), .RN(nRst), .Q(
        delta_reg[19]), .QN(n53) );
  DFC3 delta_reg_reg_17_ ( .D(delta_next[17]), .C(clk), .RN(nRst), .Q(
        delta_reg[17]), .QN(n55) );
  DFC3 delta_reg_reg_15_ ( .D(delta_next[15]), .C(clk), .RN(nRst), .Q(
        delta_reg[15]), .QN(n57) );
  DFC3 delta_reg_reg_13_ ( .D(delta_next[13]), .C(clk), .RN(nRst), .Q(
        delta_reg[13]), .QN(n59) );
  DFC3 delta_reg_reg_11_ ( .D(delta_next[11]), .C(clk), .RN(nRst), .Q(
        delta_reg[11]), .QN(n61) );
  DFC3 delta_reg_reg_9_ ( .D(delta_next[9]), .C(clk), .RN(nRst), .Q(
        delta_reg[9]), .QN(n63) );
  DFC3 delta_reg_reg_0_ ( .D(n467), .C(clk), .RN(nRst), .Q(delta_reg[0]), .QN(
        n260) );
  DFC3 state_reg_reg_1_ ( .D(n212), .C(clk), .RN(nRst), .Q(state_reg[1]), .QN(
        n38) );
  DFC3 root_reg_reg_31_ ( .D(root_next[31]), .C(clk), .RN(nRst), .Q(
        root_reg[31]) );
  DFC3 root_reg_reg_0_ ( .D(root_next[0]), .C(clk), .RN(nRst), .Q(sqroot[0])
         );
  DFC3 root_reg_reg_28_ ( .D(root_next[28]), .C(clk), .RN(nRst), .Q(
        root_reg[28]) );
  DFC3 root_reg_reg_27_ ( .D(root_next[27]), .C(clk), .RN(nRst), .Q(
        root_reg[27]) );
  DFC3 root_reg_reg_26_ ( .D(root_next[26]), .C(clk), .RN(nRst), .Q(
        root_reg[26]) );
  DFC3 root_reg_reg_25_ ( .D(n267), .C(clk), .RN(nRst), .Q(root_reg[25]) );
  DFC3 root_reg_reg_24_ ( .D(root_next[24]), .C(clk), .RN(nRst), .Q(
        root_reg[24]) );
  DFC3 root_reg_reg_23_ ( .D(n268), .C(clk), .RN(nRst), .Q(root_reg[23]) );
  DFC3 root_reg_reg_22_ ( .D(root_next[22]), .C(clk), .RN(nRst), .Q(
        root_reg[22]) );
  DFC3 root_reg_reg_21_ ( .D(root_next[21]), .C(clk), .RN(nRst), .Q(
        root_reg[21]) );
  DFC3 root_reg_reg_20_ ( .D(n242), .C(clk), .RN(nRst), .Q(root_reg[20]) );
  DFC3 root_reg_reg_19_ ( .D(n232), .C(clk), .RN(nRst), .Q(root_reg[19]) );
  DFC3 root_reg_reg_18_ ( .D(n261), .C(clk), .RN(nRst), .Q(root_reg[18]) );
  DFC3 root_reg_reg_17_ ( .D(n235), .C(clk), .RN(nRst), .Q(root_reg[17]) );
  DFC3 root_reg_reg_16_ ( .D(root_next[16]), .C(clk), .RN(nRst), .Q(sqroot[16]) );
  DFC3 root_reg_reg_14_ ( .D(root_next[14]), .C(clk), .RN(nRst), .Q(n474), 
        .QN(n233) );
  DFC3 root_reg_reg_13_ ( .D(n251), .C(clk), .RN(nRst), .Q(sqroot[13]) );
  DFC3 root_reg_reg_12_ ( .D(n250), .C(clk), .RN(nRst), .Q(n475) );
  DFC3 root_reg_reg_11_ ( .D(root_next[11]), .C(clk), .RN(nRst), .Q(sqroot[11]) );
  DFC3 root_reg_reg_10_ ( .D(root_next[10]), .C(clk), .RN(nRst), .Q(n476) );
  DFC3 root_reg_reg_9_ ( .D(n243), .C(clk), .RN(nRst), .Q(n477), .QN(n230) );
  DFC3 root_reg_reg_8_ ( .D(n241), .C(clk), .RN(nRst), .Q(n478) );
  DFC3 root_reg_reg_7_ ( .D(n252), .C(clk), .RN(nRst), .Q(sqroot[7]) );
  DFC3 root_reg_reg_6_ ( .D(n239), .C(clk), .RN(nRst), .Q(n479) );
  DFC3 root_reg_reg_5_ ( .D(n238), .C(clk), .RN(nRst), .Q(n480), .QN(n258) );
  DFC3 root_reg_reg_4_ ( .D(root_next[4]), .C(clk), .RN(nRst), .Q(n481), .QN(
        n256) );
  DFC3 root_reg_reg_3_ ( .D(root_next[3]), .C(clk), .RN(nRst), .Q(n482), .QN(
        n247) );
  DFC3 root_reg_reg_2_ ( .D(root_next[2]), .C(clk), .RN(nRst), .Q(n483) );
  DFC3 root_reg_reg_1_ ( .D(root_next[1]), .C(clk), .RN(nRst), .Q(n484) );
  DFC3 res_reg_reg_9_ ( .D(res_next[9]), .C(clk), .RN(nRst), .Q(res_reg[9]), 
        .QN(n227) );
  DFC3 res_reg_reg_8_ ( .D(res_next[8]), .C(clk), .RN(nRst), .Q(res_reg[8]) );
  DFC3 res_reg_reg_7_ ( .D(res_next[7]), .C(clk), .RN(nRst), .Q(res_reg[7]) );
  DFC3 res_reg_reg_6_ ( .D(res_next[6]), .C(clk), .RN(nRst), .Q(res_reg[6]) );
  DFC3 res_reg_reg_5_ ( .D(res_next[5]), .C(clk), .RN(nRst), .Q(res_reg[5]), 
        .QN(n249) );
  DFC3 res_reg_reg_4_ ( .D(res_next[4]), .C(clk), .RN(nRst), .Q(res_reg[4]), 
        .QN(n226) );
  DFC3 res_reg_reg_3_ ( .D(res_next[3]), .C(clk), .RN(nRst), .Q(res_reg[3]), 
        .QN(n228) );
  DFC3 res_reg_reg_30_ ( .D(res_next[30]), .C(clk), .RN(nRst), .Q(res_reg[30])
         );
  DFC3 res_reg_reg_2_ ( .D(res_next[2]), .C(clk), .RN(nRst), .Q(res_reg[2]), 
        .QN(n221) );
  DFC3 res_reg_reg_23_ ( .D(res_next[23]), .C(clk), .RN(nRst), .Q(res_reg[23])
         );
  DFC3 res_reg_reg_22_ ( .D(res_next[22]), .C(clk), .RN(nRst), .Q(res_reg[22])
         );
  DFC3 res_reg_reg_21_ ( .D(res_next[21]), .C(clk), .RN(nRst), .Q(res_reg[21])
         );
  DFC3 res_reg_reg_20_ ( .D(res_next[20]), .C(clk), .RN(nRst), .Q(res_reg[20])
         );
  DFC3 res_reg_reg_1_ ( .D(res_next[1]), .C(clk), .RN(nRst), .Q(res_reg[1]) );
  DFC3 res_reg_reg_19_ ( .D(res_next[19]), .C(clk), .RN(nRst), .Q(res_reg[19])
         );
  DFC3 res_reg_reg_18_ ( .D(res_next[18]), .C(clk), .RN(nRst), .Q(res_reg[18])
         );
  DFC3 res_reg_reg_17_ ( .D(res_next[17]), .C(clk), .RN(nRst), .Q(res_reg[17])
         );
  DFC3 res_reg_reg_16_ ( .D(res_next[16]), .C(clk), .RN(nRst), .Q(res_reg[16])
         );
  DFC3 res_reg_reg_14_ ( .D(res_next[14]), .C(clk), .RN(nRst), .Q(res_reg[14])
         );
  DFC3 res_reg_reg_13_ ( .D(res_next[13]), .C(clk), .RN(nRst), .Q(res_reg[13])
         );
  DFC3 res_reg_reg_12_ ( .D(res_next[12]), .C(clk), .RN(nRst), .Q(res_reg[12])
         );
  DFC3 res_reg_reg_11_ ( .D(res_next[11]), .C(clk), .RN(nRst), .Q(res_reg[11])
         );
  DFC3 res_reg_reg_10_ ( .D(res_next[10]), .C(clk), .RN(nRst), .Q(res_reg[10])
         );
  DFC3 res_reg_reg_0_ ( .D(res_next[0]), .C(clk), .RN(nRst), .Q(res_reg[0]) );
  DFC3 delta_reg_reg_6_ ( .D(delta_next[6]), .C(clk), .RN(nRst), .Q(
        delta_reg[6]), .QN(n66) );
  DFC3 delta_reg_reg_7_ ( .D(delta_next[7]), .C(clk), .RN(nRst), .Q(
        delta_reg[7]), .QN(n65) );
  DFC3 delta_reg_reg_5_ ( .D(n472), .C(clk), .RN(nRst), .Q(delta_reg[5]), .QN(
        n244) );
  DFC3 delta_reg_reg_4_ ( .D(n471), .C(clk), .RN(nRst), .Q(delta_reg[4]), .QN(
        n225) );
  DFC3 delta_reg_reg_3_ ( .D(n470), .C(clk), .RN(nRst), .Q(delta_reg[3]), .QN(
        n253) );
  DFC3 delta_reg_reg_2_ ( .D(n469), .C(clk), .RN(nRst), .Q(delta_reg[2]), .QN(
        n436) );
  DFC3 delta_reg_reg_1_ ( .D(n468), .C(clk), .RN(nRst), .Q(delta_reg[1]), .QN(
        n277) );
  sqroot_seq_NBITS32_DW01_inc_1 add_142 ( .A({root_reg, sqroot[16:15], n474, 
        sqroot[13:10], n477, sqroot[8:7], n215, n480, n481, n482, sqroot[2], 
        n484, sqroot[0]}), .SUM(fuo_round) );
  sqroot_seq_NBITS32_DW_cmp_5 lt_gt_109 ( .A({root_next[31:26], n267, 
        root_next[24], n268, root_next[22:21], n242, n232, n261, n235, 
        root_next[16], n246, root_next[14], n251, n250, root_next[11:10], n243, 
        n241, n252, n239, n238, root_next[4:0]}), .B({n275, res_next}), .TC(
        n_Logic0_), .GE_LT(n4), .GE_GT_EQ(n_Logic0_), .GE_LT_GT_LE(N40) );
  sqroot_seq_NBITS32_DW01_sub_5 sub_0_root_sub_0_root_sub_138 ( .A({N120, N119, 
        N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, N108, N107, 
        N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, N96, N95, N94, 
        N93, N92, N91, N90, n237}), .B({root_reg, sqroot[16:15], n474, 
        sqroot[13:10], n477, sqroot[8:7], n215, n480, n216, n482, sqroot[2:0]}), .CI(n_Logic0_), .DIFF(fuo_if_res) );
  sqroot_seq_NBITS32_DW_cmp_6 lte_110 ( .A({N73, N72, N71, N70, N69, N68, N67, 
        N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, 
        N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42}), .B({n275, 
        res_next[30:28], n264, res_next[26:0]}), .TC(n_Logic0_), .GE_LT(
        n_Logic0_), .GE_GT_EQ(n_Logic0_), .GE_LT_GT_LE(N74) );
  sqroot_seq_NBITS32_DW01_add_5 add_110 ( .A({root_next[31:26], n267, 
        root_next[24], n268, root_next[22:0]}), .B({n_Logic0_, delta_next[30], 
        n_Logic0_, delta_next[28:6], n472, n471, n470, n469, n468, n467}), 
        .CI(n_Logic0_), .SUM({N73, N72, N71, N70, N69, N68, N67, N66, N65, N64, 
        N63, N62, N61, N60, N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, 
        N49, N48, N47, N46, N45, N44, N43, N42}) );
  sqroot_seq_NBITS32_DW01_add_6 add_139 ( .A({root_reg, sqroot[16:15], n474, 
        sqroot[13:11], n476, n477, sqroot[8:7], n274, n480, n481, n482, 
        sqroot[2], n484, sqroot[0]}), .B({delta_reg[30], n_Logic0_, 
        delta_reg[28:2], n224, delta_reg[0], n_Logic0_}), .CI(n_Logic0_), 
        .SUM(fuo_if_root) );
  sqroot_seq_NBITS32_DW01_sub_7 sub_1_root_sub_0_root_sub_138 ( .A(res_reg), 
        .B({n_Logic0_, delta_reg[30], n_Logic0_, delta_reg[28:0]}), .CI(
        n_Logic0_), .DIFF({N120, N119, N118, N117, N116, N115, N114, N113, 
        N112, N111, N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, 
        N100, N99, N98, N97, N96, N95, N94, N93, N92, N91, N90, N89}) );
  DFC1 res_reg_reg_28_ ( .D(res_next[28]), .C(clk), .RN(nRst), .Q(res_reg[28])
         );
  DFC1 res_reg_reg_24_ ( .D(res_next[24]), .C(clk), .RN(nRst), .Q(res_reg[24])
         );
  DFC1 state_reg_reg_0_ ( .D(n213), .C(clk), .RN(nRst), .Q(state_reg[0]), .QN(
        n39) );
  DFC1 res_reg_reg_25_ ( .D(n245), .C(clk), .RN(nRst), .Q(res_reg[25]) );
  DFC1 res_reg_reg_26_ ( .D(res_next[26]), .C(clk), .RN(nRst), .Q(res_reg[26])
         );
  DFC1 root_reg_reg_29_ ( .D(root_next[29]), .C(clk), .RN(nRst), .Q(
        root_reg[29]) );
  DFC1 res_reg_reg_29_ ( .D(n240), .C(clk), .RN(nRst), .Q(res_reg[29]) );
  DFC1 root_reg_reg_30_ ( .D(root_next[30]), .C(clk), .RN(nRst), .Q(
        root_reg[30]) );
  DFC1 res_reg_reg_31_ ( .D(n275), .C(clk), .RN(nRst), .Q(res_reg[31]) );
  DFC3 state_reg_reg_2_ ( .D(n466), .C(clk), .RN(nRst), .Q(state_reg[2]), .QN(
        n37) );
  DFC3 res_reg_reg_27_ ( .D(n264), .C(clk), .RN(nRst), .Q(res_reg[27]) );
  DFC3 res_reg_reg_15_ ( .D(res_next[15]), .C(clk), .RN(nRst), .Q(res_reg[15])
         );
  DFC3 root_reg_reg_15_ ( .D(n246), .C(clk), .RN(nRst), .Q(n473) );
  OAI222 U264 ( .A(n4), .B(n294), .C(n45), .D(n438), .Q(delta_next[27]) );
  INV0 U265 ( .A(n273), .Q(sqroot[6]) );
  INV3 U266 ( .A(n273), .Q(n215) );
  INV6 U267 ( .A(n273), .Q(n274) );
  INV6 U268 ( .A(n479), .Q(n273) );
  NAND24 U269 ( .A(n424), .B(n423), .Q(root_next[27]) );
  INV3 U270 ( .A(n256), .Q(n216) );
  INV12 U271 ( .A(n254), .Q(sqroot[2]) );
  INV3 U272 ( .A(n262), .Q(sqroot[1]) );
  INV6 U273 ( .A(n236), .Q(n237) );
  AOI221 U274 ( .A(fuo_if_res[4]), .B(n299), .C(arg[4]), .D(n280), .Q(n361) );
  CLKIN6 U275 ( .A(n475), .Q(n217) );
  INV12 U276 ( .A(n217), .Q(sqroot[12]) );
  NAND26 U277 ( .A(n412), .B(n411), .Q(root_next[21]) );
  AOI220 U278 ( .A(fuo_if_root[0]), .B(n462), .C(sqroot[1]), .D(n291), .Q(n431) );
  NAND26 U279 ( .A(n414), .B(n413), .Q(root_next[22]) );
  NAND26 U280 ( .A(fuo_if_res[24]), .B(n299), .Q(n341) );
  BUF6 U281 ( .A(n462), .Q(n299) );
  NAND28 U282 ( .A(n347), .B(n348), .Q(n264) );
  NAND26 U283 ( .A(fuo_if_res[27]), .B(n299), .Q(n347) );
  NAND28 U284 ( .A(n324), .B(n323), .Q(res_next[16]) );
  NAND23 U285 ( .A(fuo_if_res[16]), .B(n299), .Q(n323) );
  NAND28 U286 ( .A(n356), .B(n355), .Q(res_next[30]) );
  NAND23 U287 ( .A(fuo_if_res[31]), .B(n299), .Q(n357) );
  CLKBU4 U288 ( .A(n462), .Q(n219) );
  BUF2 U289 ( .A(n462), .Q(n220) );
  INV15 U290 ( .A(n303), .Q(n462) );
  BUF6 U291 ( .A(n462), .Q(n298) );
  BUF2 U292 ( .A(n462), .Q(n266) );
  BUF2 U293 ( .A(n462), .Q(n297) );
  BUF2 U294 ( .A(n462), .Q(n300) );
  NAND23 U295 ( .A(n379), .B(n380), .Q(root_next[5]) );
  NAND24 U296 ( .A(n388), .B(n387), .Q(root_next[9]) );
  NAND23 U297 ( .A(n403), .B(n404), .Q(root_next[17]) );
  AOI221 U298 ( .A(fuo_round[19]), .B(n285), .C(root_reg[19]), .D(ready), .Q(
        n408) );
  NAND22 U299 ( .A(fuo_if_res[15]), .B(n299), .Q(n321) );
  NAND23 U300 ( .A(n358), .B(n357), .Q(n275) );
  NAND22 U301 ( .A(n312), .B(n311), .Q(res_next[10]) );
  NAND24 U302 ( .A(n398), .B(n397), .Q(root_next[14]) );
  NAND24 U303 ( .A(n418), .B(n417), .Q(root_next[24]) );
  NAND23 U304 ( .A(n426), .B(n425), .Q(root_next[28]) );
  AOI221 U305 ( .A(fuo_round[12]), .B(n284), .C(sqroot[12]), .D(n286), .Q(n394) );
  NAND23 U306 ( .A(n321), .B(n322), .Q(res_next[15]) );
  NAND23 U307 ( .A(n348), .B(n347), .Q(res_next[27]) );
  NAND26 U308 ( .A(n337), .B(n338), .Q(res_next[22]) );
  NAND26 U309 ( .A(n383), .B(n384), .Q(root_next[7]) );
  NAND26 U310 ( .A(n420), .B(n419), .Q(n267) );
  BUF8 U311 ( .A(n39), .Q(n269) );
  AOI222 U312 ( .A(fuo_if_root[11]), .B(n300), .C(sqroot[12]), .D(n291), .Q(
        n391) );
  INV3 U313 ( .A(n221), .Q(n222) );
  AOI221 U314 ( .A(n266), .B(fuo_if_root[17]), .C(n292), .D(root_reg[18]), .Q(
        n403) );
  NAND26 U315 ( .A(n409), .B(n410), .Q(root_next[20]) );
  CLKBU4 U316 ( .A(n433), .Q(n284) );
  CLKIN6 U317 ( .A(n310), .Q(n433) );
  BUF12 U318 ( .A(n433), .Q(n283) );
  INV8 U319 ( .A(n223), .Q(n224) );
  CLKIN6 U320 ( .A(n301), .Q(n302) );
  NAND23 U321 ( .A(state_reg[2]), .B(n302), .Q(n310) );
  INV3 U322 ( .A(n464), .Q(n456) );
  AOI221 U323 ( .A(fuo_round[9]), .B(n283), .C(n477), .D(n286), .Q(n388) );
  AOI221 U324 ( .A(fuo_round[17]), .B(n285), .C(root_reg[17]), .D(ready), .Q(
        n404) );
  NAND26 U325 ( .A(n405), .B(n406), .Q(root_next[18]) );
  NAND22 U326 ( .A(n430), .B(n429), .Q(root_next[30]) );
  AOI221 U327 ( .A(fuo_round[30]), .B(n284), .C(root_reg[30]), .D(ready), .Q(
        n430) );
  NAND22 U328 ( .A(n360), .B(n359), .Q(res_next[3]) );
  NAND23 U329 ( .A(n369), .B(n368), .Q(res_next[8]) );
  NAND22 U330 ( .A(n374), .B(n373), .Q(root_next[2]) );
  NAND24 U331 ( .A(n390), .B(n389), .Q(root_next[10]) );
  AOI221 U332 ( .A(fuo_round[14]), .B(n284), .C(n474), .D(n286), .Q(n398) );
  AOI221 U333 ( .A(fuo_round[23]), .B(n285), .C(root_reg[23]), .D(ready), .Q(
        n416) );
  NAND24 U334 ( .A(n422), .B(n421), .Q(root_next[26]) );
  AOI221 U335 ( .A(fuo_round[26]), .B(n284), .C(root_reg[26]), .D(ready), .Q(
        n422) );
  AOI221 U336 ( .A(fuo_round[27]), .B(n285), .C(root_reg[27]), .D(ready), .Q(
        n424) );
  AOI221 U337 ( .A(fuo_round[28]), .B(n284), .C(root_reg[28]), .D(ready), .Q(
        n426) );
  INV6 U338 ( .A(delta_reg[1]), .Q(n223) );
  CLKBU15 U339 ( .A(n452), .Q(n293) );
  AOI222 U340 ( .A(fuo_if_root[5]), .B(n220), .C(sqroot[6]), .D(n291), .Q(n379) );
  INV8 U341 ( .A(n293), .Q(n291) );
  INV6 U342 ( .A(n483), .Q(n254) );
  INV3 U343 ( .A(n228), .Q(n229) );
  OAI212 U344 ( .A(n38), .B(n456), .C(n455), .Q(n460) );
  INV3 U345 ( .A(n230), .Q(sqroot[9]) );
  BUF6 U346 ( .A(n452), .Q(n294) );
  NAND24 U347 ( .A(fuo_if_res[29]), .B(n299), .Q(n351) );
  NAND22 U348 ( .A(fuo_if_res[22]), .B(n299), .Q(n337) );
  NAND28 U349 ( .A(n330), .B(n329), .Q(res_next[19]) );
  NAND24 U350 ( .A(fuo_if_res[19]), .B(n299), .Q(n329) );
  NAND24 U351 ( .A(n376), .B(n375), .Q(root_next[3]) );
  AOI221 U352 ( .A(fuo_round[3]), .B(n283), .C(sqroot[3]), .D(n286), .Q(n376)
         );
  NAND34 U353 ( .A(n310), .B(n457), .C(n303), .Q(n454) );
  BUF2 U354 ( .A(root_next[19]), .Q(n232) );
  NAND24 U355 ( .A(n407), .B(n408), .Q(root_next[19]) );
  NAND24 U356 ( .A(N40), .B(roundup), .Q(n453) );
  INV3 U357 ( .A(n233), .Q(sqroot[14]) );
  BUF2 U358 ( .A(root_next[17]), .Q(n235) );
  NAND24 U359 ( .A(fuo_if_res[17]), .B(n299), .Q(n325) );
  CLKIN3 U360 ( .A(N89), .Q(n236) );
  NAND24 U361 ( .A(n416), .B(n415), .Q(n268) );
  NAND24 U362 ( .A(n401), .B(n402), .Q(root_next[16]) );
  AOI221 U363 ( .A(n284), .B(fuo_round[16]), .C(sqroot[16]), .D(n286), .Q(n402) );
  NAND28 U364 ( .A(n318), .B(n317), .Q(res_next[13]) );
  NAND26 U365 ( .A(fuo_if_res[13]), .B(n299), .Q(n317) );
  AOI221 U366 ( .A(fuo_if_root[29]), .B(n462), .C(root_reg[30]), .D(n291), .Q(
        n427) );
  NAND21 U367 ( .A(res_reg[0]), .B(state_reg[1]), .Q(n304) );
  BUF2 U368 ( .A(root_next[5]), .Q(n238) );
  NAND26 U369 ( .A(n393), .B(n394), .Q(root_next[12]) );
  BUF2 U370 ( .A(root_next[6]), .Q(n239) );
  BUF2 U371 ( .A(res_next[29]), .Q(n240) );
  BUF2 U372 ( .A(root_next[8]), .Q(n241) );
  BUF2 U373 ( .A(root_next[20]), .Q(n242) );
  NOR24 U374 ( .A(n279), .B(n453), .Q(n466) );
  BUF2 U375 ( .A(root_next[9]), .Q(n243) );
  NAND24 U376 ( .A(fuo_if_res[28]), .B(n299), .Q(n349) );
  NAND24 U377 ( .A(fuo_if_res[25]), .B(n299), .Q(n343) );
  NAND24 U378 ( .A(fuo_if_res[23]), .B(n299), .Q(n339) );
  AOI222 U379 ( .A(fuo_round[5]), .B(n283), .C(sqroot[5]), .D(n286), .Q(n380)
         );
  NAND26 U380 ( .A(n400), .B(n399), .Q(root_next[15]) );
  BUF2 U381 ( .A(res_next[25]), .Q(n245) );
  NAND23 U382 ( .A(fuo_if_res[12]), .B(n299), .Q(n315) );
  BUF2 U383 ( .A(root_next[15]), .Q(n246) );
  INV3 U384 ( .A(n247), .Q(sqroot[3]) );
  NAND26 U385 ( .A(fuo_if_res[18]), .B(n299), .Q(n327) );
  BUF2 U386 ( .A(root_next[12]), .Q(n250) );
  BUF2 U387 ( .A(root_next[13]), .Q(n251) );
  NAND24 U388 ( .A(n395), .B(n396), .Q(root_next[13]) );
  AOI222 U389 ( .A(fuo_round[15]), .B(n285), .C(sqroot[15]), .D(n286), .Q(n400) );
  BUF2 U390 ( .A(root_next[7]), .Q(n252) );
  NAND28 U391 ( .A(n342), .B(n341), .Q(res_next[24]) );
  NAND28 U392 ( .A(n336), .B(n335), .Q(res_next[21]) );
  AOI221 U393 ( .A(fuo_if_root[30]), .B(n462), .C(root_reg[31]), .D(n291), .Q(
        n429) );
  NAND26 U394 ( .A(n346), .B(n345), .Q(res_next[26]) );
  NAND28 U395 ( .A(n269), .B(n38), .Q(n301) );
  NAND28 U396 ( .A(n350), .B(n349), .Q(res_next[28]) );
  CLKBU15 U397 ( .A(n433), .Q(n285) );
  NAND32 U398 ( .A(state_reg[1]), .B(n269), .C(n37), .Q(n303) );
  AOI221 U399 ( .A(fuo_if_root[3]), .B(n219), .C(sqroot[4]), .D(n291), .Q(n375) );
  NAND28 U400 ( .A(n327), .B(n328), .Q(res_next[18]) );
  NAND24 U401 ( .A(fuo_if_res[21]), .B(n299), .Q(n335) );
  INV3 U402 ( .A(n256), .Q(sqroot[4]) );
  INV3 U403 ( .A(n258), .Q(sqroot[5]) );
  AOI222 U404 ( .A(fuo_if_root[9]), .B(n297), .C(sqroot[10]), .D(n291), .Q(
        n387) );
  NAND28 U405 ( .A(n351), .B(n352), .Q(res_next[29]) );
  NAND24 U406 ( .A(n378), .B(n377), .Q(root_next[4]) );
  AOI222 U407 ( .A(fuo_if_root[4]), .B(n298), .C(sqroot[5]), .D(n291), .Q(n377) );
  NAND28 U408 ( .A(n339), .B(n340), .Q(res_next[23]) );
  NAND28 U409 ( .A(n314), .B(n313), .Q(res_next[11]) );
  NAND24 U410 ( .A(fuo_if_res[11]), .B(n299), .Q(n313) );
  NAND28 U411 ( .A(n343), .B(n344), .Q(res_next[25]) );
  NAND28 U412 ( .A(n320), .B(n319), .Q(res_next[14]) );
  NAND24 U413 ( .A(fuo_if_res[14]), .B(n299), .Q(n319) );
  BUF2 U414 ( .A(root_next[18]), .Q(n261) );
  NAND26 U415 ( .A(n316), .B(n315), .Q(res_next[12]) );
  AOI212 U416 ( .A(n460), .B(n459), .C(n458), .Q(n213) );
  NAND24 U417 ( .A(fuo_if_res[20]), .B(n299), .Q(n333) );
  AOI221 U418 ( .A(fuo_round[22]), .B(n284), .C(root_reg[22]), .D(ready), .Q(
        n414) );
  AOI222 U419 ( .A(fuo_if_root[13]), .B(n220), .C(sqroot[14]), .D(n291), .Q(
        n395) );
  NAND26 U420 ( .A(n326), .B(n325), .Q(res_next[17]) );
  NAND24 U421 ( .A(n392), .B(n391), .Q(root_next[11]) );
  AOI221 U422 ( .A(fuo_round[7]), .B(n283), .C(sqroot[7]), .D(n286), .Q(n384)
         );
  NAND23 U423 ( .A(n265), .B(n302), .Q(n457) );
  CLKIN6 U424 ( .A(n484), .Q(n262) );
  AOI221 U425 ( .A(fuo_round[18]), .B(n284), .C(root_reg[18]), .D(ready), .Q(
        n406) );
  AOI222 U426 ( .A(fuo_if_root[15]), .B(n298), .C(sqroot[16]), .D(n292), .Q(
        n399) );
  AOI220 U427 ( .A(fuo_round[0]), .B(n285), .C(sqroot[0]), .D(ready), .Q(n432)
         );
  AOI221 U428 ( .A(fuo_if_root[2]), .B(n462), .C(sqroot[3]), .D(n291), .Q(n373) );
  AOI221 U429 ( .A(fuo_round[11]), .B(n285), .C(sqroot[11]), .D(n286), .Q(n392) );
  AOI221 U430 ( .A(fuo_round[10]), .B(n283), .C(sqroot[10]), .D(n286), .Q(n390) );
  AOI221 U431 ( .A(fuo_round[24]), .B(n284), .C(root_reg[24]), .D(ready), .Q(
        n418) );
  AOI221 U432 ( .A(fuo_round[4]), .B(n283), .C(sqroot[4]), .D(n286), .Q(n378)
         );
  AOI221 U433 ( .A(fuo_round[6]), .B(n283), .C(n215), .D(n286), .Q(n382) );
  AOI221 U434 ( .A(fuo_round[8]), .B(n283), .C(sqroot[8]), .D(n286), .Q(n386)
         );
  CLKBU15 U435 ( .A(n465), .Q(n286) );
  AOI221 U436 ( .A(fuo_round[20]), .B(n284), .C(root_reg[20]), .D(ready), .Q(
        n410) );
  AOI221 U437 ( .A(fuo_round[21]), .B(n285), .C(root_reg[21]), .D(ready), .Q(
        n412) );
  AOI221 U438 ( .A(fuo_round[13]), .B(n285), .C(sqroot[13]), .D(n286), .Q(n396) );
  BUF15 U439 ( .A(n465), .Q(ready) );
  CLKIN3 U440 ( .A(state_reg[2]), .Q(n265) );
  NAND22 U441 ( .A(n366), .B(n365), .Q(res_next[7]) );
  NAND22 U442 ( .A(fuo_if_res[26]), .B(n299), .Q(n345) );
  INV0 U443 ( .A(delta_next[28]), .Q(n446) );
  NAND24 U444 ( .A(n385), .B(n386), .Q(root_next[8]) );
  CLKIN3 U445 ( .A(n290), .Q(n289) );
  CLKIN3 U446 ( .A(n290), .Q(n288) );
  NAND30 U447 ( .A(n310), .B(n457), .C(n294), .Q(n367) );
  AOI220 U448 ( .A(arg[25]), .B(n282), .C(res_reg[25]), .D(n289), .Q(n344) );
  AOI220 U449 ( .A(arg[23]), .B(n282), .C(res_reg[23]), .D(n289), .Q(n340) );
  AOI220 U450 ( .A(arg[29]), .B(n282), .C(res_reg[29]), .D(n289), .Q(n352) );
  AOI220 U451 ( .A(arg[21]), .B(n282), .C(res_reg[21]), .D(n288), .Q(n336) );
  AOI220 U452 ( .A(arg[22]), .B(n281), .C(res_reg[22]), .D(n289), .Q(n338) );
  AOI220 U453 ( .A(arg[30]), .B(n282), .C(res_reg[30]), .D(n289), .Q(n356) );
  AOI220 U454 ( .A(arg[28]), .B(n281), .C(res_reg[28]), .D(n289), .Q(n350) );
  AOI220 U455 ( .A(arg[16]), .B(n282), .C(res_reg[16]), .D(n288), .Q(n324) );
  AOI220 U456 ( .A(arg[18]), .B(n282), .C(res_reg[18]), .D(n288), .Q(n328) );
  AOI220 U457 ( .A(arg[26]), .B(n281), .C(res_reg[26]), .D(n289), .Q(n346) );
  AOI220 U458 ( .A(arg[20]), .B(n281), .C(res_reg[20]), .D(n288), .Q(n334) );
  AOI220 U459 ( .A(arg[31]), .B(n281), .C(res_reg[31]), .D(n289), .Q(n358) );
  NOR40 U460 ( .A(n451), .B(n450), .C(n449), .D(n448), .Q(n464) );
  CLKIN3 U461 ( .A(n293), .Q(n292) );
  BUF2 U462 ( .A(n461), .Q(n280) );
  BUF2 U463 ( .A(n461), .Q(n282) );
  BUF2 U464 ( .A(n461), .Q(n281) );
  INV3 U465 ( .A(n367), .Q(n290) );
  NAND41 U466 ( .A(n442), .B(n441), .C(n440), .D(n439), .Q(n451) );
  NOR40 U467 ( .A(delta_next[6]), .B(delta_next[7]), .C(n472), .D(n471), .Q(
        n441) );
  NOR40 U468 ( .A(delta_next[15]), .B(delta_next[14]), .C(delta_next[13]), .D(
        delta_next[12]), .Q(n439) );
  NOR40 U469 ( .A(delta_next[11]), .B(delta_next[10]), .C(delta_next[9]), .D(
        delta_next[8]), .Q(n440) );
  BUF2 U470 ( .A(n452), .Q(n295) );
  BUF2 U471 ( .A(n452), .Q(n296) );
  NOR40 U472 ( .A(delta_next[23]), .B(delta_next[22]), .C(delta_next[21]), .D(
        delta_next[20]), .Q(n443) );
  NOR40 U473 ( .A(delta_next[27]), .B(delta_next[26]), .C(delta_next[25]), .D(
        delta_next[24]), .Q(n447) );
  NOR40 U474 ( .A(delta_next[19]), .B(delta_next[18]), .C(delta_next[17]), .D(
        delta_next[16]), .Q(n444) );
  INV3 U475 ( .A(n437), .Q(n461) );
  AOI220 U476 ( .A(arg[12]), .B(n280), .C(res_reg[12]), .D(n288), .Q(n316) );
  AOI220 U477 ( .A(arg[2]), .B(n281), .C(n222), .D(n289), .Q(n354) );
  AOI220 U478 ( .A(fuo_round[29]), .B(n285), .C(root_reg[29]), .D(ready), .Q(
        n428) );
  AOI220 U479 ( .A(fuo_round[31]), .B(n284), .C(root_reg[31]), .D(ready), .Q(
        n435) );
  NAND22 U480 ( .A(n372), .B(n371), .Q(root_next[1]) );
  AOI220 U481 ( .A(arg[11]), .B(n280), .C(res_reg[11]), .D(n288), .Q(n314) );
  AOI220 U482 ( .A(arg[19]), .B(n281), .C(res_reg[19]), .D(n288), .Q(n330) );
  AOI220 U483 ( .A(arg[24]), .B(n281), .C(res_reg[24]), .D(n289), .Q(n342) );
  AOI220 U484 ( .A(arg[15]), .B(n280), .C(res_reg[15]), .D(n288), .Q(n322) );
  AOI220 U485 ( .A(arg[14]), .B(n280), .C(res_reg[14]), .D(n288), .Q(n320) );
  NAND24 U486 ( .A(n381), .B(n382), .Q(root_next[6]) );
  AOI220 U487 ( .A(arg[13]), .B(n280), .C(res_reg[13]), .D(n288), .Q(n318) );
  AOI220 U488 ( .A(arg[27]), .B(n282), .C(res_reg[27]), .D(n289), .Q(n348) );
  AOI220 U489 ( .A(fuo_if_res[5]), .B(n462), .C(arg[5]), .D(n280), .Q(n362) );
  AOI220 U490 ( .A(arg[1]), .B(n282), .C(res_reg[1]), .D(n288), .Q(n332) );
  AOI220 U491 ( .A(arg[17]), .B(n281), .C(res_reg[17]), .D(n288), .Q(n326) );
  AOI220 U492 ( .A(arg[8]), .B(n281), .C(res_reg[8]), .D(n289), .Q(n369) );
  AOI220 U493 ( .A(arg[6]), .B(n281), .C(res_reg[6]), .D(n289), .Q(n364) );
  AOI220 U494 ( .A(arg[7]), .B(n282), .C(res_reg[7]), .D(n289), .Q(n366) );
  AOI220 U495 ( .A(arg[3]), .B(n282), .C(n229), .D(n289), .Q(n360) );
  AOI220 U496 ( .A(arg[10]), .B(n280), .C(res_reg[10]), .D(n288), .Q(n312) );
  AOI220 U497 ( .A(arg[0]), .B(n280), .C(fuo_if_res[0]), .D(n300), .Q(n309) );
  AOI220 U498 ( .A(n265), .B(n307), .C(res_reg[0]), .D(n283), .Q(n308) );
  OAI311 U499 ( .A(n464), .B(state_reg[2]), .C(n38), .D(n463), .Q(n212) );
  NOR20 U500 ( .A(n299), .B(n280), .Q(n463) );
  LOGIC0 U501 ( .Q(n_Logic0_) );
  LOGIC1 U502 ( .Q(n4) );
  AOI222 U503 ( .A(fuo_if_root[10]), .B(n266), .C(sqroot[11]), .D(n291), .Q(
        n389) );
  AOI222 U504 ( .A(fuo_if_root[24]), .B(n462), .C(root_reg[25]), .D(n292), .Q(
        n417) );
  AOI222 U505 ( .A(fuo_if_root[6]), .B(n266), .C(sqroot[7]), .D(n291), .Q(n381) );
  NOR40 U506 ( .A(n470), .B(n469), .C(n467), .D(n468), .Q(n442) );
  CLKIN6 U507 ( .A(n478), .Q(n270) );
  INV12 U508 ( .A(n270), .Q(sqroot[8]) );
  CLKBU15 U509 ( .A(n473), .Q(sqroot[15]) );
  CLKBU15 U510 ( .A(n476), .Q(sqroot[10]) );
  AOI222 U511 ( .A(fuo_if_root[7]), .B(n297), .C(sqroot[8]), .D(n291), .Q(n383) );
  NAND31 U512 ( .A(state_reg[0]), .B(n38), .C(n265), .Q(n437) );
  CLKIN1 U513 ( .A(n269), .Q(n459) );
  NAND20 U514 ( .A(res_reg[0]), .B(n269), .Q(n306) );
  NOR21 U515 ( .A(n294), .B(n456), .Q(n278) );
  INV3 U516 ( .A(n278), .Q(n279) );
  NAND28 U517 ( .A(n333), .B(n334), .Q(res_next[20]) );
  INV3 U518 ( .A(N74), .Q(n455) );
  AOI220 U519 ( .A(fuo_round[1]), .B(n283), .C(sqroot[1]), .D(n286), .Q(n372)
         );
  AOI220 U520 ( .A(fuo_round[2]), .B(n283), .C(sqroot[2]), .D(n286), .Q(n374)
         );
  AOI220 U521 ( .A(fuo_if_root[1]), .B(n462), .C(sqroot[2]), .D(n291), .Q(n371) );
  INV15 U522 ( .A(n454), .Q(n438) );
  INV6 U523 ( .A(n457), .Q(n465) );
  NAND33 U524 ( .A(state_reg[0]), .B(state_reg[1]), .C(n265), .Q(n452) );
  OAI222 U525 ( .A(n294), .B(n253), .C(n438), .D(n277), .Q(n468) );
  OAI222 U526 ( .A(n296), .B(n225), .C(n438), .D(n436), .Q(n469) );
  OAI222 U527 ( .A(n296), .B(n244), .C(n438), .D(n253), .Q(n470) );
  OAI222 U528 ( .A(n296), .B(n66), .C(n438), .D(n225), .Q(n471) );
  OAI222 U529 ( .A(n296), .B(n65), .C(n438), .D(n244), .Q(n472) );
  OAI222 U530 ( .A(n63), .B(n296), .C(n65), .D(n438), .Q(delta_next[7]) );
  OAI222 U531 ( .A(n64), .B(n296), .C(n66), .D(n438), .Q(delta_next[6]) );
  CLKIN3 U532 ( .A(state_reg[0]), .Q(n305) );
  OAI222 U533 ( .A(state_reg[1]), .B(n306), .C(n305), .D(n304), .Q(n307) );
  NAND22 U534 ( .A(n309), .B(n308), .Q(res_next[0]) );
  NAND22 U535 ( .A(fuo_if_res[10]), .B(n299), .Q(n311) );
  NAND22 U536 ( .A(fuo_if_res[1]), .B(n462), .Q(n331) );
  NAND22 U537 ( .A(n332), .B(n331), .Q(res_next[1]) );
  NAND22 U538 ( .A(fuo_if_res[2]), .B(n299), .Q(n353) );
  NAND22 U539 ( .A(n354), .B(n353), .Q(res_next[2]) );
  NAND22 U540 ( .A(fuo_if_res[30]), .B(n299), .Q(n355) );
  NAND22 U541 ( .A(fuo_if_res[3]), .B(n462), .Q(n359) );
  OAI212 U542 ( .A(n290), .B(n226), .C(n361), .Q(res_next[4]) );
  OAI212 U543 ( .A(n290), .B(n249), .C(n362), .Q(res_next[5]) );
  NAND22 U544 ( .A(fuo_if_res[6]), .B(n299), .Q(n363) );
  NAND22 U545 ( .A(n364), .B(n363), .Q(res_next[6]) );
  NAND22 U546 ( .A(fuo_if_res[7]), .B(n299), .Q(n365) );
  NAND22 U547 ( .A(fuo_if_res[8]), .B(n299), .Q(n368) );
  AOI222 U548 ( .A(fuo_if_res[9]), .B(n299), .C(arg[9]), .D(n280), .Q(n370) );
  OAI212 U549 ( .A(n290), .B(n227), .C(n370), .Q(res_next[9]) );
  AOI222 U550 ( .A(fuo_if_root[8]), .B(n300), .C(sqroot[9]), .D(n291), .Q(n385) );
  AOI222 U551 ( .A(fuo_if_root[12]), .B(n266), .C(sqroot[13]), .D(n291), .Q(
        n393) );
  AOI222 U552 ( .A(fuo_if_root[14]), .B(n300), .C(sqroot[15]), .D(n292), .Q(
        n397) );
  AOI222 U553 ( .A(fuo_if_root[16]), .B(n297), .C(root_reg[17]), .D(n292), .Q(
        n401) );
  AOI222 U554 ( .A(fuo_if_root[18]), .B(n297), .C(root_reg[19]), .D(n292), .Q(
        n405) );
  AOI222 U555 ( .A(fuo_if_root[19]), .B(n462), .C(root_reg[20]), .D(n292), .Q(
        n407) );
  AOI222 U556 ( .A(fuo_if_root[20]), .B(n462), .C(root_reg[21]), .D(n292), .Q(
        n409) );
  AOI222 U557 ( .A(fuo_if_root[21]), .B(n462), .C(root_reg[22]), .D(n292), .Q(
        n411) );
  AOI222 U558 ( .A(fuo_if_root[22]), .B(n219), .C(root_reg[23]), .D(n292), .Q(
        n413) );
  AOI222 U559 ( .A(fuo_if_root[23]), .B(n462), .C(root_reg[24]), .D(n292), .Q(
        n415) );
  AOI222 U560 ( .A(fuo_round[25]), .B(n285), .C(root_reg[25]), .D(ready), .Q(
        n420) );
  AOI222 U561 ( .A(fuo_if_root[25]), .B(n462), .C(root_reg[26]), .D(n292), .Q(
        n419) );
  AOI222 U562 ( .A(fuo_if_root[26]), .B(n462), .C(root_reg[27]), .D(n292), .Q(
        n421) );
  AOI222 U563 ( .A(fuo_if_root[27]), .B(n462), .C(root_reg[28]), .D(n292), .Q(
        n423) );
  AOI222 U564 ( .A(fuo_if_root[28]), .B(n462), .C(root_reg[29]), .D(n292), .Q(
        n425) );
  NAND22 U565 ( .A(n428), .B(n427), .Q(root_next[29]) );
  NAND22 U566 ( .A(n432), .B(n431), .Q(root_next[0]) );
  NAND22 U567 ( .A(fuo_if_root[31]), .B(n299), .Q(n434) );
  NAND22 U568 ( .A(n435), .B(n434), .Q(root_next[31]) );
  OAI222 U569 ( .A(n438), .B(n260), .C(n294), .D(n436), .Q(n467) );
  OAI222 U570 ( .A(n62), .B(n296), .C(n64), .D(n438), .Q(delta_next[8]) );
  OAI222 U571 ( .A(n61), .B(n296), .C(n63), .D(n438), .Q(delta_next[9]) );
  OAI222 U572 ( .A(n60), .B(n294), .C(n62), .D(n438), .Q(delta_next[10]) );
  OAI222 U573 ( .A(n59), .B(n295), .C(n61), .D(n438), .Q(delta_next[11]) );
  OAI222 U574 ( .A(n58), .B(n294), .C(n60), .D(n438), .Q(delta_next[12]) );
  OAI222 U575 ( .A(n57), .B(n294), .C(n59), .D(n438), .Q(delta_next[13]) );
  OAI222 U576 ( .A(n56), .B(n295), .C(n58), .D(n438), .Q(delta_next[14]) );
  OAI222 U577 ( .A(n55), .B(n295), .C(n57), .D(n438), .Q(delta_next[15]) );
  OAI222 U578 ( .A(n54), .B(n295), .C(n56), .D(n438), .Q(delta_next[16]) );
  OAI222 U579 ( .A(n53), .B(n295), .C(n55), .D(n438), .Q(delta_next[17]) );
  OAI222 U580 ( .A(n52), .B(n295), .C(n54), .D(n438), .Q(delta_next[18]) );
  OAI222 U581 ( .A(n51), .B(n295), .C(n53), .D(n438), .Q(delta_next[19]) );
  OAI222 U582 ( .A(n50), .B(n295), .C(n52), .D(n438), .Q(delta_next[20]) );
  OAI222 U583 ( .A(n49), .B(n295), .C(n51), .D(n438), .Q(delta_next[21]) );
  OAI222 U584 ( .A(n48), .B(n295), .C(n50), .D(n438), .Q(delta_next[22]) );
  OAI222 U585 ( .A(n47), .B(n295), .C(n49), .D(n438), .Q(delta_next[23]) );
  OAI222 U586 ( .A(n46), .B(n294), .C(n48), .D(n438), .Q(delta_next[24]) );
  OAI222 U587 ( .A(n45), .B(n294), .C(n47), .D(n438), .Q(delta_next[25]) );
  OAI222 U588 ( .A(n44), .B(n294), .C(n46), .D(n438), .Q(delta_next[26]) );
  OAI222 U589 ( .A(n42), .B(n294), .C(n44), .D(n438), .Q(delta_next[28]) );
  OAI212 U590 ( .A(n42), .B(n438), .C(n437), .Q(delta_next[30]) );
  NAND22 U591 ( .A(n444), .B(n443), .Q(n450) );
  CLKIN3 U592 ( .A(delta_next[30]), .Q(n445) );
  NAND22 U593 ( .A(n446), .B(n445), .Q(n449) );
  CLKIN3 U594 ( .A(n447), .Q(n448) );
  OAI212 U595 ( .A(start), .B(n457), .C(n37), .Q(n458) );
endmodule

