
module sqroot_comb_NBITS16_DW01_inc_6 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;
  wire   n1, n2, n3, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n21, n23, n24, n25, n28, n29, n33;

  CLKIN0 U47 ( .A(A[3]), .Q(n23) );
  NAND20 U48 ( .A(A[0]), .B(n18), .Q(n17) );
  NAND21 U49 ( .A(A[0]), .B(n10), .Q(n9) );
  NAND22 U50 ( .A(A[0]), .B(n15), .Q(n14) );
  NAND21 U51 ( .A(A[0]), .B(n25), .Q(n24) );
  NAND21 U52 ( .A(A[0]), .B(n7), .Q(n6) );
  CLKIN3 U53 ( .A(A[2]), .Q(n28) );
  XNR21 U54 ( .A(A[7]), .B(n6), .Q(SUM[7]) );
  CLKIN0 U55 ( .A(n18), .Q(n19) );
  NOR20 U56 ( .A(n28), .B(n33), .Q(n25) );
  INV0 U57 ( .A(n11), .Q(n10) );
  INV2 U58 ( .A(n3), .Q(n2) );
  NAND20 U59 ( .A(n7), .B(A[7]), .Q(n3) );
  INV0 U60 ( .A(A[6]), .Q(n8) );
  INV2 U61 ( .A(n1), .Q(SUM[8]) );
  NOR21 U62 ( .A(n16), .B(n19), .Q(n15) );
  NOR21 U63 ( .A(n21), .B(n33), .Q(n18) );
  INV0 U64 ( .A(A[4]), .Q(n16) );
  NOR21 U65 ( .A(n8), .B(n11), .Q(n7) );
  CLKIN0 U66 ( .A(A[1]), .Q(n33) );
  NAND22 U67 ( .A(n18), .B(n12), .Q(n11) );
  NOR21 U68 ( .A(n13), .B(n16), .Q(n12) );
  XOR21 U69 ( .A(n28), .B(n29), .Q(SUM[2]) );
  NAND20 U70 ( .A(A[0]), .B(A[1]), .Q(n29) );
  XOR21 U71 ( .A(n13), .B(n14), .Q(SUM[5]) );
  XNR20 U72 ( .A(n33), .B(A[0]), .Q(SUM[1]) );
  XOR21 U73 ( .A(n8), .B(n9), .Q(SUM[6]) );
  XOR21 U74 ( .A(n23), .B(n24), .Q(SUM[3]) );
  XOR21 U75 ( .A(n16), .B(n17), .Q(SUM[4]) );
  INV0 U76 ( .A(A[5]), .Q(n13) );
  NAND20 U77 ( .A(A[0]), .B(n2), .Q(n1) );
  NAND20 U78 ( .A(A[2]), .B(A[3]), .Q(n21) );
endmodule


module sqroot_comb_NBITS16 ( arg, roundup, sqroot );
  input [15:0] arg;
  output [8:0] sqroot;
  input roundup;
  wire   N711, N712, N713, N714, N715, N716, N717, N718, lt_gt_52_A_7_,
         lt_gt_52_A_4_, lt_gt_52_A_1_, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1472,
         SYNOPSYS_UNCONNECTED_1;

  sqroot_comb_NBITS16_DW01_inc_6 add_53 ( .A({n1472, n908, n878, n879, n887, 
        n888, n1470, n718, n712}), .SUM({N718, N717, N716, N715, N714, N713, 
        N712, N711, SYNOPSYS_UNCONNECTED_1}) );
  INV3 U643 ( .A(n1097), .Q(n755) );
  NAND33 U644 ( .A(n1148), .B(n746), .C(n1149), .Q(n1096) );
  INV10 U645 ( .A(n1179), .Q(n759) );
  INV4 U646 ( .A(n954), .Q(n970) );
  NAND26 U647 ( .A(n951), .B(n950), .Q(n954) );
  INV10 U648 ( .A(n706), .Q(n1104) );
  NAND23 U649 ( .A(n1280), .B(n851), .Q(n1288) );
  BUF6 U650 ( .A(n1273), .Q(n851) );
  INV12 U651 ( .A(n1135), .Q(n1169) );
  CLKIN6 U652 ( .A(n1354), .Q(n1337) );
  NAND24 U653 ( .A(n1000), .B(n1009), .Q(n1023) );
  NAND33 U654 ( .A(n1110), .B(n1109), .C(n1137), .Q(n1124) );
  INV3 U655 ( .A(n654), .Q(n651) );
  NAND24 U656 ( .A(n1279), .B(n1278), .Q(n1313) );
  NAND32 U657 ( .A(n1231), .B(n1230), .C(n887), .Q(n1278) );
  INV6 U658 ( .A(n1111), .Q(n731) );
  CLKIN10 U659 ( .A(n1228), .Q(n1240) );
  NAND42 U660 ( .A(n1012), .B(n988), .C(n987), .D(n756), .Q(n625) );
  INV3 U661 ( .A(n684), .Q(n1400) );
  INV6 U662 ( .A(n1448), .Q(n626) );
  INV6 U663 ( .A(arg[13]), .Q(n855) );
  CLKBU12 U664 ( .A(n949), .Q(n909) );
  NAND23 U665 ( .A(n800), .B(n910), .Q(n1445) );
  INV4 U666 ( .A(n1445), .Q(n836) );
  NAND22 U667 ( .A(n1445), .B(n837), .Q(n838) );
  INV12 U668 ( .A(n1469), .Q(n1448) );
  INV10 U669 ( .A(n1412), .Q(n789) );
  NAND24 U670 ( .A(n1039), .B(n1036), .Q(n1051) );
  NAND22 U671 ( .A(n1118), .B(n627), .Q(n628) );
  NAND22 U672 ( .A(n1117), .B(n1116), .Q(n629) );
  NAND24 U673 ( .A(n628), .B(n629), .Q(n769) );
  CLKIN6 U674 ( .A(n1116), .Q(n627) );
  XNR22 U675 ( .A(lt_gt_52_A_7_), .B(n1048), .Q(n669) );
  NOR24 U676 ( .A(n630), .B(arg[13]), .Q(n631) );
  NOR23 U677 ( .A(n631), .B(n914), .Q(n917) );
  INV8 U678 ( .A(arg[12]), .Q(n630) );
  NOR32 U679 ( .A(arg[12]), .B(arg[10]), .C(arg[11]), .Q(n914) );
  CLKIN12 U680 ( .A(n1180), .Q(n1097) );
  INV8 U681 ( .A(n1007), .Q(n1005) );
  CLKIN6 U682 ( .A(n1171), .Q(n632) );
  CLKIN15 U683 ( .A(n1155), .Q(n1171) );
  BUF6 U684 ( .A(n1155), .Q(n728) );
  NAND26 U685 ( .A(n1034), .B(n1035), .Q(n1038) );
  NAND24 U686 ( .A(n1034), .B(n1027), .Q(n1039) );
  NAND33 U687 ( .A(n1150), .B(n755), .C(n1179), .Q(n1188) );
  INV15 U688 ( .A(arg[13]), .Q(n856) );
  NAND23 U689 ( .A(n871), .B(n912), .Q(n913) );
  INV12 U690 ( .A(n1469), .Q(n949) );
  NAND33 U691 ( .A(n934), .B(n935), .C(n1469), .Q(n940) );
  OAI2112 U692 ( .A(arg[12]), .B(arg[13]), .C(arg[14]), .D(arg[15]), .Q(n912)
         );
  INV6 U693 ( .A(n1108), .Q(n633) );
  CLKIN6 U694 ( .A(n1108), .Q(n1120) );
  NAND28 U695 ( .A(n863), .B(n1106), .Q(n1108) );
  INV4 U696 ( .A(n1134), .Q(n1132) );
  NAND28 U697 ( .A(n1114), .B(n1115), .Q(n1134) );
  NAND24 U698 ( .A(n641), .B(n642), .Q(n1260) );
  NAND28 U699 ( .A(arg[12]), .B(arg[15]), .Q(n927) );
  INV12 U700 ( .A(n663), .Q(n1416) );
  NAND23 U701 ( .A(n1311), .B(n908), .Q(n771) );
  INV4 U702 ( .A(n625), .Q(n994) );
  NAND28 U703 ( .A(n1021), .B(n999), .Q(n1010) );
  INV3 U704 ( .A(n661), .Q(n634) );
  INV6 U705 ( .A(n853), .Q(n661) );
  NAND26 U706 ( .A(n716), .B(n888), .Q(n1377) );
  NAND34 U707 ( .A(n1038), .B(n1059), .C(lt_gt_52_A_4_), .Q(n1074) );
  CLKIN15 U708 ( .A(arg[10]), .Q(n864) );
  INV4 U709 ( .A(n1067), .Q(n783) );
  CLKIN3 U710 ( .A(n1384), .Q(n635) );
  INV12 U711 ( .A(n1384), .Q(n1264) );
  NAND22 U712 ( .A(n636), .B(n637), .Q(n638) );
  NAND24 U713 ( .A(n638), .B(n915), .Q(n916) );
  INV3 U714 ( .A(arg[14]), .Q(n636) );
  INV3 U715 ( .A(arg[15]), .Q(n637) );
  INV8 U716 ( .A(n1038), .Q(n1061) );
  NOR32 U717 ( .A(n1260), .B(n853), .C(n1261), .Q(n1266) );
  CLKIN3 U718 ( .A(n1168), .Q(n1160) );
  NAND23 U719 ( .A(n1197), .B(n1160), .Q(n1161) );
  CLKIN15 U720 ( .A(n1419), .Q(n1057) );
  CLKIN6 U721 ( .A(n1419), .Q(n888) );
  INV4 U722 ( .A(n1098), .Q(n1189) );
  NAND26 U723 ( .A(n760), .B(n1098), .Q(n1093) );
  NAND23 U724 ( .A(n666), .B(n667), .Q(n1049) );
  IMUX24 U725 ( .A(n877), .B(n1136), .S(n1470), .Q(n1133) );
  INV6 U726 ( .A(n1169), .Q(n773) );
  NAND23 U727 ( .A(n652), .B(n653), .Q(n1223) );
  INV15 U728 ( .A(n1421), .Q(lt_gt_52_A_1_) );
  INV4 U729 ( .A(n1234), .Q(n1140) );
  INV6 U730 ( .A(n1404), .Q(n1396) );
  INV4 U731 ( .A(lt_gt_52_A_1_), .Q(n750) );
  INV3 U732 ( .A(n1421), .Q(n857) );
  NAND23 U733 ( .A(n1162), .B(n1161), .Q(n1163) );
  OAI212 U734 ( .A(n1133), .B(n827), .C(n1270), .Q(n683) );
  NAND24 U735 ( .A(n1108), .B(arg[6]), .Q(n1110) );
  NAND23 U736 ( .A(n835), .B(n799), .Q(n800) );
  NAND26 U737 ( .A(n745), .B(n878), .Q(n748) );
  CLKIN4 U738 ( .A(n1055), .Q(n745) );
  INV12 U739 ( .A(n1029), .Q(n818) );
  INV12 U740 ( .A(n1070), .Q(n1064) );
  INV10 U741 ( .A(n832), .Q(n762) );
  CLKIN2 U742 ( .A(n1064), .Q(n817) );
  CLKIN3 U743 ( .A(n1228), .Q(n713) );
  INV2 U744 ( .A(n1097), .Q(n687) );
  NOR32 U745 ( .A(n689), .B(n1368), .C(n1367), .Q(n882) );
  NAND21 U746 ( .A(n1258), .B(n1259), .Q(n641) );
  NAND24 U747 ( .A(n639), .B(n640), .Q(n642) );
  INV1 U748 ( .A(n1258), .Q(n639) );
  INV4 U749 ( .A(n1259), .Q(n640) );
  CLKIN8 U750 ( .A(n884), .Q(n886) );
  INV6 U751 ( .A(n1237), .Q(n1225) );
  NAND22 U752 ( .A(n650), .B(n654), .Q(n653) );
  NAND24 U753 ( .A(n1394), .B(n889), .Q(n1374) );
  INV2 U754 ( .A(n1033), .Q(n1072) );
  INV2 U755 ( .A(n1013), .Q(n1004) );
  CLKIN15 U756 ( .A(n835), .Q(n861) );
  INV12 U757 ( .A(n1256), .Q(n853) );
  CLKIN6 U758 ( .A(n1057), .Q(n828) );
  NAND34 U759 ( .A(n1294), .B(n1293), .C(n908), .Q(n1287) );
  NAND24 U760 ( .A(n769), .B(n824), .Q(n1216) );
  CLKIN8 U761 ( .A(n769), .Q(n1270) );
  NAND28 U762 ( .A(n822), .B(n1157), .Q(n1166) );
  INV4 U763 ( .A(n1154), .Q(n722) );
  NAND23 U764 ( .A(n1470), .B(n1192), .Q(n1332) );
  NAND22 U765 ( .A(n1019), .B(n1016), .Q(n847) );
  CLKBU15 U766 ( .A(n1216), .Q(n905) );
  NAND23 U767 ( .A(n1421), .B(n1241), .Q(n715) );
  INV6 U768 ( .A(n1190), .Q(n1308) );
  NAND24 U769 ( .A(n1301), .B(n1302), .Q(n1147) );
  INV6 U770 ( .A(n1274), .Q(n1277) );
  INV1 U771 ( .A(n1059), .Q(n1060) );
  INV1 U772 ( .A(n1173), .Q(n1181) );
  INV6 U773 ( .A(n847), .Q(n848) );
  OAI212 U774 ( .A(n1137), .B(n877), .C(n1124), .Q(n1126) );
  INV12 U775 ( .A(n1467), .Q(n1466) );
  NOR23 U776 ( .A(n795), .B(n880), .Q(n881) );
  INV6 U777 ( .A(n992), .Q(n997) );
  INV3 U778 ( .A(n646), .Q(n1100) );
  NOR23 U779 ( .A(arg[14]), .B(arg[13]), .Q(n741) );
  NAND22 U780 ( .A(n1055), .B(n746), .Q(n747) );
  NOR23 U781 ( .A(n986), .B(n881), .Q(n987) );
  NAND23 U782 ( .A(n989), .B(n910), .Q(n990) );
  NAND24 U783 ( .A(n918), .B(n1017), .Q(n1008) );
  NOR21 U784 ( .A(n962), .B(arg[11]), .Q(n701) );
  NAND26 U785 ( .A(n976), .B(n975), .Q(n1101) );
  NAND24 U786 ( .A(n971), .B(n884), .Q(n976) );
  INV6 U787 ( .A(arg[8]), .Q(n1017) );
  BUF8 U788 ( .A(n1101), .Q(n757) );
  INV3 U789 ( .A(n1073), .Q(n1077) );
  NAND23 U790 ( .A(n1181), .B(n878), .Q(n1198) );
  NAND26 U791 ( .A(n1338), .B(n1377), .Q(n1339) );
  NAND24 U792 ( .A(n1146), .B(n737), .Q(n1302) );
  NAND24 U793 ( .A(n835), .B(n797), .Q(n1383) );
  NAND21 U794 ( .A(n824), .B(n1345), .Q(n797) );
  INV3 U795 ( .A(n682), .Q(n648) );
  NAND24 U796 ( .A(n1470), .B(n1413), .Q(n1388) );
  NAND22 U797 ( .A(n1252), .B(n859), .Q(n1255) );
  INV3 U798 ( .A(n1329), .Q(n1298) );
  INV3 U799 ( .A(n823), .Q(n824) );
  INV6 U800 ( .A(n1442), .Q(n1395) );
  INV0 U801 ( .A(n1345), .Q(n808) );
  INV10 U802 ( .A(n1385), .Q(n1345) );
  CLKIN12 U803 ( .A(n716), .Q(n1394) );
  INV15 U804 ( .A(n911), .Q(n878) );
  BUF15 U805 ( .A(n1403), .Q(n911) );
  INV10 U806 ( .A(n1036), .Q(n1058) );
  NAND21 U807 ( .A(n1447), .B(n803), .Q(n1457) );
  OAI210 U808 ( .A(n1061), .B(n1060), .C(n737), .Q(n1062) );
  CLKIN1 U809 ( .A(n1466), .Q(n862) );
  OAI212 U810 ( .A(n1346), .B(n1345), .C(n699), .Q(n643) );
  CLKIN4 U811 ( .A(n778), .Q(n738) );
  INV6 U812 ( .A(arg[15]), .Q(n644) );
  BUF15 U813 ( .A(n949), .Q(n910) );
  NAND23 U814 ( .A(n1040), .B(n649), .Q(n1052) );
  INV3 U815 ( .A(arg[15]), .Q(n1172) );
  NAND24 U816 ( .A(n646), .B(n1018), .Q(n1065) );
  CLKBU15 U817 ( .A(n941), .Q(n854) );
  INV10 U818 ( .A(n955), .Q(n941) );
  NAND26 U819 ( .A(n1154), .B(n1171), .Q(n1157) );
  CLKIN10 U820 ( .A(n1156), .Q(n1154) );
  NAND24 U821 ( .A(n1448), .B(n777), .Q(n950) );
  INV2 U822 ( .A(n1032), .Q(n1043) );
  INV3 U823 ( .A(n1020), .Q(n993) );
  NAND23 U824 ( .A(n1028), .B(n983), .Q(n988) );
  INV6 U825 ( .A(n1402), .Q(n756) );
  NAND24 U826 ( .A(n732), .B(n733), .Q(n1112) );
  CLKIN10 U827 ( .A(n1402), .Q(n884) );
  INV6 U828 ( .A(n885), .Q(n887) );
  INV2 U829 ( .A(n1009), .Q(n1011) );
  CLKIN6 U830 ( .A(n1010), .Q(n736) );
  NAND28 U831 ( .A(n1404), .B(n694), .Q(n663) );
  CLKIN2 U832 ( .A(n888), .Q(n860) );
  NAND24 U833 ( .A(n1440), .B(n811), .Q(n1458) );
  INV3 U834 ( .A(n1068), .Q(n907) );
  NAND22 U835 ( .A(n1062), .B(n649), .Q(n1068) );
  NAND28 U836 ( .A(n1069), .B(n1022), .Q(n1082) );
  NAND23 U837 ( .A(n1246), .B(arg[3]), .Q(n845) );
  INV2 U838 ( .A(n739), .Q(n740) );
  INV8 U839 ( .A(n1178), .Q(n1150) );
  BUF2 U840 ( .A(n861), .Q(n645) );
  CLKIN6 U841 ( .A(n1142), .Q(n827) );
  NAND26 U842 ( .A(n783), .B(n906), .Q(n784) );
  INV12 U843 ( .A(n753), .Q(n1454) );
  CLKIN6 U844 ( .A(n1282), .Q(n656) );
  AOI212 U845 ( .A(n886), .B(arg[8]), .C(n1081), .Q(n646) );
  INV12 U846 ( .A(n1271), .Q(n901) );
  INV4 U847 ( .A(n1293), .Q(n1292) );
  INV3 U848 ( .A(n1052), .Q(n1041) );
  OAI311 U849 ( .A(n1183), .B(n1450), .C(n1182), .D(n1198), .Q(n1186) );
  CLKIN3 U850 ( .A(n1244), .Q(n1245) );
  NAND28 U851 ( .A(n1166), .B(n823), .Q(n1193) );
  BUF2 U852 ( .A(n1296), .Q(n647) );
  IMUX24 U853 ( .A(n1382), .B(n1383), .S(n648), .Q(n1387) );
  NAND32 U854 ( .A(n1038), .B(n1059), .C(n887), .Q(n649) );
  CLKIN3 U855 ( .A(n719), .Q(n699) );
  INV8 U856 ( .A(n1065), .Q(n1069) );
  NAND23 U857 ( .A(n1184), .B(n1188), .Q(n1185) );
  NAND28 U858 ( .A(n1283), .B(n718), .Q(n752) );
  NAND26 U859 ( .A(n763), .B(n764), .Q(n1056) );
  NAND28 U860 ( .A(n758), .B(n759), .Q(n760) );
  NAND24 U861 ( .A(n674), .B(n675), .Q(n677) );
  INV3 U862 ( .A(n1317), .Q(n674) );
  NAND24 U863 ( .A(n651), .B(n1147), .Q(n652) );
  INV3 U864 ( .A(n1147), .Q(n650) );
  NAND28 U865 ( .A(n1112), .B(n1124), .Q(n1151) );
  NAND26 U866 ( .A(n1159), .B(n737), .Q(n1168) );
  INV4 U867 ( .A(n939), .Q(n974) );
  NAND23 U868 ( .A(n1243), .B(n1362), .Q(n1328) );
  NAND24 U869 ( .A(n1008), .B(n991), .Q(n992) );
  NAND26 U870 ( .A(n767), .B(n1374), .Q(n1341) );
  INV6 U871 ( .A(n1350), .Q(n1353) );
  INV10 U872 ( .A(n892), .Q(n1156) );
  INV6 U873 ( .A(n1313), .Q(n1315) );
  XOR22 U874 ( .A(n1291), .B(n879), .Q(n654) );
  NAND22 U875 ( .A(n807), .B(n1282), .Q(n657) );
  NAND28 U876 ( .A(n656), .B(n655), .Q(n658) );
  NAND28 U877 ( .A(n657), .B(n658), .Q(n1283) );
  CLKIN6 U878 ( .A(n807), .Q(n655) );
  NAND24 U879 ( .A(n937), .B(n730), .Q(n659) );
  NAND33 U880 ( .A(n924), .B(n939), .C(n660), .Q(n729) );
  INV6 U881 ( .A(n659), .Q(n660) );
  INV3 U882 ( .A(n1450), .Q(n730) );
  NAND23 U883 ( .A(n923), .B(n922), .Q(n924) );
  CLKIN3 U884 ( .A(n1317), .Q(n1290) );
  NAND28 U885 ( .A(n672), .B(n673), .Q(n1442) );
  NAND23 U886 ( .A(n1044), .B(n809), .Q(n1045) );
  NAND23 U887 ( .A(n1217), .B(n1218), .Q(n1219) );
  NAND28 U888 ( .A(n835), .B(n678), .Q(n1412) );
  NAND28 U889 ( .A(n1057), .B(n1056), .Q(n1092) );
  NAND26 U890 ( .A(n1290), .B(n878), .Q(n1314) );
  NAND28 U891 ( .A(n1037), .B(n1058), .Q(n1032) );
  INV6 U892 ( .A(n1039), .Q(n1037) );
  INV4 U893 ( .A(n958), .Q(n934) );
  INV4 U894 ( .A(n940), .Q(n953) );
  NAND21 U895 ( .A(n1469), .B(n991), .Q(n980) );
  INV2 U896 ( .A(n626), .Q(n823) );
  NAND28 U897 ( .A(n933), .B(n964), .Q(n1469) );
  INV4 U898 ( .A(n1417), .Q(n1459) );
  CLKIN12 U899 ( .A(n1286), .Q(n1273) );
  OAI222 U900 ( .A(n909), .B(n985), .C(arg[10]), .D(n984), .Q(n986) );
  CLKIN3 U901 ( .A(n1301), .Q(n815) );
  XNR22 U902 ( .A(n909), .B(n1385), .Q(n1380) );
  NAND24 U903 ( .A(n1284), .B(n786), .Q(n1294) );
  NAND23 U904 ( .A(n1269), .B(n1271), .Q(n1230) );
  NAND22 U905 ( .A(n1194), .B(n1193), .Q(n1196) );
  NAND34 U906 ( .A(n1263), .B(n910), .C(n1262), .Q(n1384) );
  XNR22 U907 ( .A(n813), .B(n980), .Q(n1012) );
  OAI221 U908 ( .A(n1469), .B(n957), .C(arg[10]), .D(n997), .Q(n960) );
  XNR21 U909 ( .A(n1008), .B(n626), .Q(n977) );
  NOR20 U910 ( .A(n878), .B(n626), .Q(n794) );
  CLKIN12 U911 ( .A(n824), .Q(n979) );
  NAND26 U912 ( .A(n1373), .B(n1372), .Q(n1379) );
  INV6 U913 ( .A(n796), .Q(n787) );
  BUF2 U914 ( .A(n1012), .Q(n692) );
  INV2 U915 ( .A(n1362), .Q(n1364) );
  NAND22 U916 ( .A(n982), .B(n878), .Q(n985) );
  INV3 U917 ( .A(arg[10]), .Q(n991) );
  NAND22 U918 ( .A(n1054), .B(n762), .Q(n763) );
  CLKIN3 U919 ( .A(n701), .Q(n957) );
  INV6 U920 ( .A(n1006), .Q(n890) );
  INV3 U921 ( .A(n1318), .Q(n1325) );
  NAND26 U922 ( .A(n861), .B(arg[0]), .Q(n1423) );
  NAND33 U923 ( .A(n1015), .B(n848), .C(n711), .Q(n1106) );
  NAND24 U924 ( .A(n742), .B(n1429), .Q(n744) );
  CLKIN6 U925 ( .A(n861), .Q(n662) );
  NAND26 U926 ( .A(n1071), .B(n817), .Q(n1102) );
  INV2 U927 ( .A(n910), .Q(n879) );
  NAND24 U928 ( .A(n1355), .B(n686), .Q(n1370) );
  NOR22 U929 ( .A(n801), .B(n1453), .Q(n1461) );
  INV2 U930 ( .A(n861), .Q(n712) );
  XOR31 U931 ( .A(n911), .B(n1173), .C(n1163), .Q(n1164) );
  NAND28 U932 ( .A(n747), .B(n748), .Q(n832) );
  INV2 U933 ( .A(n1010), .Q(n1024) );
  INV12 U934 ( .A(n757), .Q(n711) );
  NOR21 U935 ( .A(n1370), .B(n883), .Q(n1371) );
  XOR22 U936 ( .A(n645), .B(n1456), .Q(sqroot[0]) );
  NAND28 U937 ( .A(n1344), .B(n1343), .Q(n1385) );
  INV2 U938 ( .A(n1322), .Q(n796) );
  AOI312 U939 ( .A(n1409), .B(n896), .C(n662), .D(n1408), .Q(n1415) );
  CLKIN12 U940 ( .A(n905), .Q(n703) );
  NAND24 U941 ( .A(lt_gt_52_A_1_), .B(n1470), .Q(n1259) );
  INV0 U942 ( .A(n1413), .Q(n788) );
  INV3 U943 ( .A(n1388), .Q(n1390) );
  CLKIN6 U944 ( .A(n1339), .Q(n1342) );
  NAND24 U945 ( .A(n798), .B(n1341), .Q(n1343) );
  NAND24 U946 ( .A(n877), .B(n773), .Q(n774) );
  NAND20 U947 ( .A(n1209), .B(n888), .Q(n1212) );
  NAND28 U948 ( .A(n818), .B(n819), .Q(n821) );
  NAND22 U949 ( .A(n1047), .B(n665), .Q(n666) );
  NAND22 U950 ( .A(n664), .B(n669), .Q(n667) );
  INV4 U951 ( .A(n1047), .Q(n664) );
  INV3 U952 ( .A(n669), .Q(n665) );
  NAND24 U953 ( .A(n1067), .B(n907), .Q(n785) );
  INV6 U954 ( .A(n750), .Q(n718) );
  INV4 U955 ( .A(n1434), .Q(n742) );
  INV3 U956 ( .A(n683), .Q(n1275) );
  INV12 U957 ( .A(n1413), .Q(n1247) );
  INV6 U958 ( .A(n1423), .Q(n1422) );
  NAND28 U959 ( .A(n751), .B(n752), .Q(n753) );
  CLKIN2 U960 ( .A(n1444), .Q(n749) );
  CLKIN6 U961 ( .A(n1424), .Q(n1425) );
  INV12 U962 ( .A(n1269), .Q(n1142) );
  NOR24 U963 ( .A(n875), .B(n861), .Q(n1431) );
  NAND28 U964 ( .A(n1444), .B(lt_gt_52_A_4_), .Q(n1338) );
  CLKIN6 U965 ( .A(n1405), .Q(n1444) );
  CLKIN12 U966 ( .A(n1193), .Q(n1175) );
  INV6 U967 ( .A(n695), .Q(n668) );
  INV12 U968 ( .A(n1270), .Q(n695) );
  NAND26 U969 ( .A(n1422), .B(n895), .Q(n1426) );
  NAND22 U970 ( .A(n808), .B(n719), .Q(n1386) );
  NAND26 U971 ( .A(n1169), .B(n1137), .Q(n1144) );
  NOR23 U972 ( .A(n889), .B(n1224), .Q(n781) );
  INV12 U973 ( .A(n1144), .Q(n1224) );
  OAI210 U974 ( .A(n888), .B(n1210), .C(arg[4]), .Q(n1211) );
  NAND24 U975 ( .A(n1311), .B(n1450), .Q(n1329) );
  INV15 U976 ( .A(n776), .Q(n1271) );
  NOR22 U977 ( .A(arg[15]), .B(arg[14]), .Q(n873) );
  INV15 U978 ( .A(arg[15]), .Q(n866) );
  NAND28 U979 ( .A(n714), .B(n715), .Q(n716) );
  NAND26 U980 ( .A(n828), .B(n829), .Q(n830) );
  NAND26 U981 ( .A(n1405), .B(n737), .Q(n1256) );
  NAND24 U982 ( .A(n806), .B(n1299), .Q(n1310) );
  OAI212 U983 ( .A(n647), .B(n1295), .C(n1294), .Q(n1331) );
  NAND22 U984 ( .A(n1434), .B(n1435), .Q(n743) );
  NAND28 U985 ( .A(n1387), .B(n1386), .Q(n1404) );
  NAND24 U986 ( .A(n743), .B(n744), .Q(n1436) );
  NAND23 U987 ( .A(n1412), .B(n1413), .Q(n790) );
  INV2 U988 ( .A(n1179), .Q(n1202) );
  NAND22 U989 ( .A(n1393), .B(n1394), .Q(n672) );
  NAND26 U990 ( .A(n670), .B(n671), .Q(n673) );
  CLKIN6 U991 ( .A(n1393), .Q(n670) );
  CLKIN3 U992 ( .A(n1394), .Q(n671) );
  NAND21 U993 ( .A(n1317), .B(n878), .Q(n676) );
  NAND24 U994 ( .A(n676), .B(n677), .Q(n807) );
  INV0 U995 ( .A(n878), .Q(n675) );
  NAND26 U996 ( .A(n1289), .B(n1288), .Q(n1317) );
  INV2 U997 ( .A(n1348), .Q(n1351) );
  OAI222 U998 ( .A(n662), .B(n1407), .C(n896), .D(n1407), .Q(n1408) );
  NAND30 U999 ( .A(n835), .B(n1358), .C(roundup), .Q(n801) );
  NAND20 U1000 ( .A(n835), .B(n1430), .Q(n1428) );
  NAND23 U1001 ( .A(n835), .B(n1392), .Q(n1393) );
  CLKIN4 U1002 ( .A(n680), .Q(n825) );
  NAND22 U1003 ( .A(n1418), .B(n888), .Q(n1414) );
  CLKIN15 U1004 ( .A(n890), .Q(n891) );
  NAND26 U1005 ( .A(n1420), .B(n860), .Q(n1441) );
  CLKIN12 U1006 ( .A(n1143), .Q(n1141) );
  INV2 U1007 ( .A(n1377), .Q(n1375) );
  NAND23 U1008 ( .A(n1303), .B(n1314), .Q(n1304) );
  OAI211 U1009 ( .A(n1316), .B(n1315), .C(n1314), .Q(n690) );
  NAND24 U1010 ( .A(n1073), .B(n793), .Q(n1149) );
  BUF2 U1011 ( .A(n635), .Q(n719) );
  CLKIN6 U1012 ( .A(n884), .Q(n885) );
  CLKIN6 U1013 ( .A(lt_gt_52_A_4_), .Q(n737) );
  NAND28 U1014 ( .A(n790), .B(n791), .Q(n1418) );
  NAND28 U1015 ( .A(n789), .B(n788), .Q(n791) );
  NAND24 U1016 ( .A(n826), .B(n1081), .Q(n1059) );
  NAND24 U1017 ( .A(n1353), .B(n878), .Q(n1362) );
  NAND26 U1018 ( .A(n680), .B(n1244), .Q(n1421) );
  BUF6 U1019 ( .A(n1411), .Q(n678) );
  CLKIN6 U1020 ( .A(n1205), .Q(n679) );
  CLKIN12 U1021 ( .A(n679), .Q(n680) );
  INV10 U1022 ( .A(n978), .Q(n1029) );
  INV6 U1023 ( .A(n906), .Q(n707) );
  INV3 U1024 ( .A(n826), .Q(n906) );
  NAND24 U1025 ( .A(n1142), .B(n901), .Q(n1231) );
  OAI222 U1026 ( .A(n885), .B(n1017), .C(n979), .D(n1033), .Q(n1016) );
  NAND23 U1027 ( .A(n1033), .B(n909), .Q(n1019) );
  NAND34 U1028 ( .A(n1005), .B(n891), .C(n977), .Q(n978) );
  NAND28 U1029 ( .A(n1049), .B(n830), .Q(n1098) );
  CLKIN6 U1030 ( .A(n1285), .Q(n1322) );
  INV4 U1031 ( .A(n1230), .Q(n1146) );
  INV1 U1032 ( .A(n878), .Q(n746) );
  INV3 U1033 ( .A(n1028), .Q(n819) );
  INV3 U1034 ( .A(arg[7]), .Q(n1087) );
  INV3 U1035 ( .A(n1371), .Q(n1460) );
  XOR22 U1036 ( .A(n749), .B(n800), .Q(n681) );
  INV0 U1037 ( .A(n1454), .Q(n1358) );
  INV3 U1038 ( .A(n937), .Q(n972) );
  INV6 U1039 ( .A(lt_gt_52_A_7_), .Q(n1450) );
  BUF2 U1040 ( .A(n1381), .Q(n682) );
  NAND21 U1041 ( .A(n1263), .B(n1262), .Q(n1381) );
  BUF2 U1042 ( .A(n1361), .Q(n869) );
  NAND23 U1043 ( .A(n1381), .B(n824), .Q(n1361) );
  XOR22 U1044 ( .A(n1391), .B(n860), .Q(n1392) );
  INV2 U1045 ( .A(n921), .Q(n880) );
  INV1 U1046 ( .A(n1361), .Q(n1346) );
  NAND24 U1047 ( .A(n1281), .B(n1280), .Q(n1291) );
  NAND23 U1048 ( .A(n1228), .B(n901), .Q(n1262) );
  BUF15 U1049 ( .A(n799), .Q(n896) );
  NAND24 U1050 ( .A(n1098), .B(n1099), .Q(n1128) );
  XNR22 U1051 ( .A(n1432), .B(n1431), .Q(n1438) );
  NAND34 U1052 ( .A(n1015), .B(n848), .C(n711), .Q(n706) );
  NAND22 U1053 ( .A(n749), .B(n824), .Q(n1406) );
  NOR33 U1054 ( .A(n861), .B(n702), .C(n1347), .Q(n1398) );
  NAND24 U1055 ( .A(n1423), .B(n720), .Q(n1424) );
  OAI312 U1056 ( .A(n873), .B(n1398), .C(n1399), .D(n1397), .Q(n684) );
  AOI222 U1057 ( .A(n803), .B(n1447), .C(n1459), .D(n1458), .Q(n1464) );
  OAI212 U1058 ( .A(n883), .B(n1370), .C(roundup), .Q(n1463) );
  NOR22 U1059 ( .A(n1379), .B(n1380), .Q(n1382) );
  NOR23 U1060 ( .A(n1210), .B(n867), .Q(n831) );
  NAND26 U1061 ( .A(n731), .B(arg[7]), .Q(n733) );
  OAI221 U1062 ( .A(n849), .B(n1457), .C(n1449), .D(n1465), .Q(n1455) );
  INV0 U1063 ( .A(n1400), .Q(n849) );
  AOI212 U1064 ( .A(n997), .B(n956), .C(n1448), .Q(n961) );
  NAND24 U1065 ( .A(n663), .B(n1441), .Q(n810) );
  AOI211 U1066 ( .A(n1236), .B(n1235), .C(n724), .Q(n1238) );
  CLKIN3 U1067 ( .A(n1241), .Q(n1236) );
  NAND34 U1068 ( .A(n1142), .B(n901), .C(n695), .Q(n1280) );
  CLKIN3 U1069 ( .A(n1339), .Q(n798) );
  CLKIN6 U1070 ( .A(n1389), .Q(n685) );
  INV6 U1071 ( .A(n1410), .Q(n1389) );
  NAND24 U1072 ( .A(n1267), .B(n1268), .Q(n1327) );
  XOR31 U1073 ( .A(n860), .B(n1237), .C(n850), .Q(n1226) );
  NAND28 U1074 ( .A(n1247), .B(n898), .Q(n767) );
  INV0 U1075 ( .A(n1337), .Q(n686) );
  INV1 U1076 ( .A(n1188), .Q(n1182) );
  INV1 U1077 ( .A(n1138), .Q(n868) );
  OAI2112 U1078 ( .A(n824), .B(n632), .C(n1096), .D(n1090), .Q(n688) );
  CLKIN0 U1079 ( .A(n910), .Q(n802) );
  INV6 U1080 ( .A(n1107), .Q(n1105) );
  NAND22 U1081 ( .A(n717), .B(n746), .Q(n1174) );
  CLKIN6 U1082 ( .A(n1174), .Q(n1195) );
  OAI210 U1083 ( .A(n895), .B(n1310), .C(n1309), .Q(n689) );
  NAND21 U1084 ( .A(n958), .B(n873), .Q(n959) );
  CLKIN2 U1085 ( .A(n1185), .Q(n1200) );
  INV3 U1086 ( .A(n924), .Q(n973) );
  INV1 U1087 ( .A(n1159), .Q(n1113) );
  INV0 U1088 ( .A(n1273), .Q(n691) );
  CLKIN6 U1089 ( .A(n1057), .Q(n693) );
  INV3 U1090 ( .A(n878), .Q(n694) );
  NOR21 U1091 ( .A(n740), .B(n1102), .Q(n1103) );
  CLKIN0 U1092 ( .A(n1332), .Q(n1333) );
  NAND28 U1093 ( .A(n1222), .B(n1221), .Q(n1244) );
  NOR42 U1094 ( .A(n709), .B(n1036), .C(n707), .D(n1050), .Q(n1031) );
  NOR23 U1095 ( .A(n876), .B(n868), .Q(n867) );
  XOR31 U1096 ( .A(n737), .B(n1152), .C(n1113), .Q(n1117) );
  INV0 U1097 ( .A(n1152), .Q(n1125) );
  NOR22 U1098 ( .A(n1322), .B(n758), .Q(n696) );
  NAND28 U1099 ( .A(n725), .B(n726), .Q(n1036) );
  NAND22 U1100 ( .A(n1028), .B(n1029), .Q(n725) );
  XNR22 U1101 ( .A(arg[8]), .B(n1402), .Q(n826) );
  INV6 U1102 ( .A(n1102), .Q(n1022) );
  INV6 U1103 ( .A(n1443), .Q(n799) );
  BUF2 U1104 ( .A(n1291), .Q(n768) );
  NOR21 U1105 ( .A(n749), .B(n824), .Q(n697) );
  BUF2 U1106 ( .A(n1433), .Q(n698) );
  AOI212 U1107 ( .A(n1351), .B(n878), .C(n723), .Q(n1352) );
  NAND24 U1108 ( .A(n1051), .B(n1032), .Q(n1055) );
  INV3 U1109 ( .A(n1146), .Q(n700) );
  NAND24 U1110 ( .A(n1024), .B(n1023), .Q(n1050) );
  CLKIN3 U1111 ( .A(n966), .Q(n841) );
  NAND23 U1112 ( .A(n841), .B(n840), .Q(n843) );
  INV3 U1113 ( .A(n962), .Q(n963) );
  CLKIN15 U1114 ( .A(arg[11]), .Q(n981) );
  INV0 U1115 ( .A(n1353), .Q(n702) );
  INV2 U1116 ( .A(n1359), .Q(n1360) );
  XOR31 U1117 ( .A(n824), .B(n1166), .C(n1194), .Q(n1170) );
  CLKIN6 U1118 ( .A(n1217), .Q(n1296) );
  INV0 U1119 ( .A(n1140), .Q(n724) );
  INV4 U1120 ( .A(n1023), .Q(n1001) );
  INV3 U1121 ( .A(n1012), .Q(n1000) );
  NOR33 U1122 ( .A(n901), .B(lt_gt_52_A_4_), .C(n703), .Q(n704) );
  NOR24 U1123 ( .A(n1215), .B(n704), .Q(n1222) );
  INV2 U1124 ( .A(n1184), .Q(n1183) );
  INV1 U1125 ( .A(n1053), .Q(n705) );
  NAND24 U1126 ( .A(n1313), .B(n1312), .Q(n1282) );
  INV6 U1127 ( .A(n1075), .Q(n1053) );
  CLKIN0 U1128 ( .A(n1225), .Q(n708) );
  INV2 U1129 ( .A(n1027), .Q(n709) );
  XOR22 U1130 ( .A(n878), .B(n643), .Q(n1347) );
  CLKIN0 U1131 ( .A(n1072), .Q(n792) );
  INV6 U1132 ( .A(n1178), .Q(n754) );
  CLKIN3 U1133 ( .A(n994), .Q(n710) );
  OAI222 U1134 ( .A(n1089), .B(n693), .C(n1057), .D(n1088), .Q(n1090) );
  CLKIN15 U1135 ( .A(n1379), .Q(n835) );
  NAND21 U1136 ( .A(n1317), .B(n694), .Q(n1319) );
  INV2 U1137 ( .A(n1101), .Q(n1018) );
  OAI210 U1138 ( .A(arg[7]), .B(n1122), .C(n885), .Q(n1078) );
  NOR24 U1139 ( .A(n698), .B(n861), .Q(n1434) );
  INV1 U1140 ( .A(n1372), .Q(n723) );
  NAND21 U1141 ( .A(n691), .B(n750), .Q(n751) );
  INV6 U1142 ( .A(n1130), .Q(n1138) );
  NOR42 U1143 ( .A(n860), .B(n1394), .C(n1264), .D(n853), .Q(n1242) );
  NAND24 U1144 ( .A(n857), .B(n1248), .Q(n714) );
  INV3 U1145 ( .A(n1239), .Q(n1248) );
  OAI211 U1146 ( .A(n755), .B(n1150), .C(n1177), .Q(n717) );
  NAND28 U1147 ( .A(n1148), .B(n1149), .Q(n1180) );
  NAND21 U1148 ( .A(n633), .B(n1119), .Q(n1121) );
  NAND23 U1149 ( .A(n1419), .B(n1004), .Q(n1091) );
  XOR31 U1150 ( .A(n909), .B(n1074), .C(n1053), .Q(n1076) );
  INV0 U1151 ( .A(n895), .Q(n720) );
  INV2 U1152 ( .A(lt_gt_52_A_1_), .Q(n895) );
  NAND26 U1153 ( .A(n1138), .B(n1134), .Q(n1135) );
  INV4 U1154 ( .A(n1054), .Q(n761) );
  NAND21 U1155 ( .A(n940), .B(n936), .Q(n937) );
  INV6 U1156 ( .A(n1063), .Q(n1071) );
  BUF2 U1157 ( .A(n1111), .Q(n902) );
  CLKBU15 U1158 ( .A(n1050), .Q(n721) );
  INV6 U1159 ( .A(n1128), .Q(n1114) );
  CLKIN6 U1160 ( .A(n1030), .Q(n1027) );
  NAND28 U1161 ( .A(n774), .B(n775), .Q(n776) );
  NAND24 U1162 ( .A(n819), .B(n818), .Q(n726) );
  OAI312 U1163 ( .A(n1325), .B(n852), .C(n1324), .D(n1323), .Q(n727) );
  INV6 U1164 ( .A(n729), .Q(n971) );
  OAI211 U1165 ( .A(n1470), .B(n1238), .C(n708), .Q(n1239) );
  NAND24 U1166 ( .A(n1201), .B(n1470), .Q(n1217) );
  NAND33 U1167 ( .A(n1009), .B(n1450), .C(n1000), .Q(n1020) );
  NAND21 U1168 ( .A(n1188), .B(n1189), .Q(n1307) );
  NAND28 U1169 ( .A(n820), .B(n821), .Q(n1013) );
  NAND22 U1170 ( .A(n1029), .B(n1028), .Q(n820) );
  XNR22 U1171 ( .A(arg[4]), .B(n1470), .Q(n1241) );
  INV12 U1172 ( .A(n1437), .Q(n1470) );
  NAND22 U1173 ( .A(n1111), .B(n1087), .Q(n732) );
  NAND28 U1174 ( .A(n1013), .B(n694), .Q(n1070) );
  INV3 U1175 ( .A(n1051), .Q(n1042) );
  NAND21 U1176 ( .A(n1134), .B(n1206), .Q(n876) );
  CLKIN6 U1177 ( .A(n948), .Q(n777) );
  NOR21 U1178 ( .A(arg[10]), .B(n813), .Q(n734) );
  NOR23 U1179 ( .A(n735), .B(n949), .Q(n812) );
  INV3 U1180 ( .A(n734), .Q(n735) );
  INV3 U1181 ( .A(arg[11]), .Q(n813) );
  NAND28 U1182 ( .A(n633), .B(n1082), .Q(n1419) );
  NAND23 U1183 ( .A(n1167), .B(n1168), .Q(n1176) );
  INV6 U1184 ( .A(n947), .Q(n778) );
  NAND23 U1185 ( .A(n1151), .B(n1154), .Q(n1159) );
  NOR21 U1186 ( .A(n1100), .B(n757), .Q(n739) );
  OAI211 U1187 ( .A(n1127), .B(n1128), .C(n1206), .Q(n1129) );
  NOR33 U1188 ( .A(n996), .B(n812), .C(n995), .Q(n920) );
  INV6 U1189 ( .A(n919), .Q(n995) );
  NAND23 U1190 ( .A(n681), .B(n824), .Q(n803) );
  NAND34 U1191 ( .A(n822), .B(n1157), .C(n879), .Q(n1197) );
  INV6 U1192 ( .A(n1150), .Q(n822) );
  NAND24 U1193 ( .A(n761), .B(n832), .Q(n764) );
  INV3 U1194 ( .A(n1167), .Q(n1158) );
  NOR23 U1195 ( .A(n834), .B(n1306), .Q(n1309) );
  CLKIN6 U1196 ( .A(n1176), .Q(n1194) );
  NAND24 U1197 ( .A(n1115), .B(n1114), .Q(n1139) );
  NAND28 U1198 ( .A(n1156), .B(n1155), .Q(n1178) );
  NOR24 U1199 ( .A(n893), .B(n872), .Q(n1116) );
  AOI212 U1200 ( .A(n1032), .B(n721), .C(n1031), .Q(n1048) );
  INV6 U1201 ( .A(n765), .Q(n766) );
  OAI212 U1202 ( .A(arg[0]), .B(n861), .C(arg[1]), .Q(n1427) );
  NAND34 U1203 ( .A(n1071), .B(n817), .C(n1069), .Q(n1119) );
  CLKIN3 U1204 ( .A(lt_gt_52_A_1_), .Q(n852) );
  NOR32 U1205 ( .A(n1065), .B(n1064), .C(n1063), .Q(n1066) );
  INV3 U1206 ( .A(n908), .Q(n758) );
  XOR22 U1207 ( .A(n1277), .B(n1232), .Q(n1233) );
  NAND24 U1208 ( .A(n1233), .B(n713), .Q(n1263) );
  NOR33 U1209 ( .A(arg[6]), .B(n1105), .C(n1104), .Q(n765) );
  NOR24 U1210 ( .A(n766), .B(n1103), .Q(n1111) );
  NAND28 U1211 ( .A(n845), .B(n846), .Q(n1413) );
  NAND28 U1212 ( .A(n844), .B(n1257), .Q(n846) );
  NAND28 U1213 ( .A(n770), .B(n1450), .Q(n772) );
  NAND28 U1214 ( .A(n771), .B(n772), .Q(n1318) );
  CLKIN6 U1215 ( .A(n1311), .Q(n770) );
  NAND24 U1216 ( .A(n1136), .B(n1169), .Q(n775) );
  NAND24 U1217 ( .A(n1294), .B(n1293), .Q(n1311) );
  AOI212 U1218 ( .A(n1126), .B(n860), .C(n1125), .Q(n1136) );
  CLKIN12 U1219 ( .A(n1418), .Q(n1420) );
  NAND26 U1220 ( .A(n836), .B(n697), .Q(n839) );
  INV3 U1221 ( .A(n882), .Q(n883) );
  NAND21 U1222 ( .A(n948), .B(n778), .Q(n779) );
  NAND22 U1223 ( .A(n777), .B(n738), .Q(n780) );
  NAND22 U1224 ( .A(n779), .B(n780), .Q(n951) );
  NOR32 U1225 ( .A(n1142), .B(n782), .C(n1141), .Q(n1145) );
  INV3 U1226 ( .A(n781), .Q(n782) );
  INV0 U1227 ( .A(n888), .Q(n889) );
  NAND28 U1228 ( .A(n784), .B(n785), .Q(n1155) );
  NAND43 U1229 ( .A(n661), .B(n767), .C(n1254), .D(n1255), .Q(n1268) );
  NOR24 U1230 ( .A(n787), .B(n851), .Q(n786) );
  INV2 U1231 ( .A(n1331), .Q(n1297) );
  INV2 U1232 ( .A(n792), .Q(n793) );
  INV3 U1233 ( .A(n794), .Q(n795) );
  NAND24 U1234 ( .A(n838), .B(n839), .Q(n1446) );
  CLKIN6 U1235 ( .A(n1272), .Q(n1289) );
  NOR33 U1236 ( .A(n909), .B(n1275), .C(n1284), .Q(n1276) );
  XOR31 U1237 ( .A(lt_gt_52_A_7_), .B(n1185), .C(n1199), .Q(n1201) );
  OAI222 U1238 ( .A(n887), .B(n1230), .C(n1231), .D(lt_gt_52_A_4_), .Q(n1229)
         );
  NAND22 U1239 ( .A(n804), .B(n805), .Q(n806) );
  INV0 U1240 ( .A(n1300), .Q(n804) );
  INV2 U1241 ( .A(n1330), .Q(n805) );
  INV6 U1242 ( .A(n1246), .Q(n844) );
  NAND23 U1243 ( .A(n949), .B(n981), .Q(n919) );
  OAI222 U1244 ( .A(n1350), .B(n635), .C(n694), .D(n1264), .Q(n1254) );
  NAND23 U1245 ( .A(n1138), .B(n1134), .Q(n1437) );
  OAI212 U1246 ( .A(n1264), .B(n1338), .C(n1361), .Q(n1265) );
  NAND28 U1247 ( .A(n1005), .B(n891), .Q(n1402) );
  NAND26 U1248 ( .A(n1005), .B(n891), .Q(n1026) );
  INV6 U1249 ( .A(n913), .Q(n933) );
  NAND22 U1250 ( .A(n855), .B(n945), .Q(n943) );
  NOR33 U1251 ( .A(n825), .B(arg[2]), .C(n1245), .Q(n1246) );
  NAND24 U1252 ( .A(arg[12]), .B(n925), .Q(n926) );
  NAND26 U1253 ( .A(n1289), .B(n787), .Q(n1293) );
  NAND22 U1254 ( .A(n746), .B(n1036), .Q(n809) );
  INV6 U1255 ( .A(n810), .Q(n811) );
  OAI222 U1256 ( .A(n1352), .B(n1353), .C(n1359), .D(n1351), .Q(n1399) );
  XNR22 U1257 ( .A(n1017), .B(n1026), .Q(n1034) );
  INV0 U1258 ( .A(n1406), .Q(n1409) );
  INV8 U1259 ( .A(arg[12]), .Q(n945) );
  OAI311 U1260 ( .A(n1007), .B(arg[8]), .C(n890), .D(arg[9]), .Q(n1025) );
  INV15 U1261 ( .A(arg[15]), .Q(n814) );
  INV3 U1262 ( .A(n815), .Q(n816) );
  CLKIN3 U1263 ( .A(n989), .Q(n1028) );
  OAI220 U1264 ( .A(arg[4]), .B(n1212), .C(n1437), .D(n1211), .Q(n1213) );
  NAND21 U1265 ( .A(n1350), .B(n694), .Q(n1359) );
  XNR20 U1266 ( .A(n1410), .B(n1470), .Q(n1411) );
  CLKIN3 U1267 ( .A(n1470), .Q(n898) );
  NAND21 U1268 ( .A(n1470), .B(n1257), .Q(n1258) );
  NAND21 U1269 ( .A(n1202), .B(n1135), .Q(n1218) );
  NAND22 U1270 ( .A(n690), .B(n1319), .Q(n1324) );
  INV6 U1271 ( .A(n990), .Q(n998) );
  NAND24 U1272 ( .A(n1077), .B(n1076), .Q(n1148) );
  AOI212 U1273 ( .A(arg[11]), .B(n910), .C(n911), .Q(n938) );
  OAI2112 U1274 ( .A(n879), .B(n681), .C(n663), .D(n1395), .Q(n1401) );
  AOI312 U1275 ( .A(n1302), .B(n1312), .C(n816), .D(n1300), .Q(n1303) );
  IMUX22 U1276 ( .A(n1365), .B(n1366), .S(n1451), .Q(n1367) );
  AOI222 U1277 ( .A(n787), .B(n852), .C(n1321), .D(n718), .Q(n1323) );
  BUF2 U1278 ( .A(n903), .Q(n850) );
  OAI222 U1279 ( .A(n1186), .B(n1187), .C(n908), .D(n1200), .Q(n1190) );
  NAND21 U1280 ( .A(n878), .B(n1051), .Q(n1046) );
  INV6 U1281 ( .A(n1139), .Q(n872) );
  INV0 U1282 ( .A(n721), .Q(n829) );
  NAND34 U1283 ( .A(n1140), .B(n1207), .C(arg[5]), .Q(n1143) );
  CLKIN6 U1284 ( .A(n867), .Q(n1207) );
  NAND20 U1285 ( .A(n1454), .B(n908), .Q(n1365) );
  NAND20 U1286 ( .A(n1454), .B(n1450), .Q(n1366) );
  NOR31 U1287 ( .A(n833), .B(n1191), .C(n898), .Q(n834) );
  INV0 U1288 ( .A(n1308), .Q(n833) );
  INV6 U1289 ( .A(n1349), .Q(n1372) );
  OAI212 U1290 ( .A(n1399), .B(n1398), .C(n1450), .Q(n1355) );
  INV1 U1291 ( .A(n697), .Q(n837) );
  INV6 U1292 ( .A(n1151), .Q(n1153) );
  AOI312 U1293 ( .A(n685), .B(n1388), .C(n1377), .D(n1376), .Q(n1378) );
  NAND22 U1294 ( .A(n967), .B(n966), .Q(n842) );
  NAND24 U1295 ( .A(n842), .B(n843), .Q(n968) );
  INV3 U1296 ( .A(n967), .Q(n840) );
  NOR23 U1297 ( .A(n866), .B(arg[14]), .Q(n865) );
  NAND32 U1298 ( .A(n865), .B(n870), .C(n855), .Q(n871) );
  XNR22 U1299 ( .A(arg[10]), .B(n949), .Q(n921) );
  XNR20 U1300 ( .A(arg[2]), .B(n718), .Q(n1435) );
  NAND21 U1301 ( .A(lt_gt_52_A_1_), .B(n1331), .Q(n1334) );
  XNR22 U1302 ( .A(n887), .B(n1378), .Q(n1443) );
  NAND22 U1303 ( .A(n1330), .B(n1329), .Q(n1336) );
  NOR33 U1304 ( .A(n1335), .B(n1298), .C(n1297), .Q(n1299) );
  AOI222 U1305 ( .A(arg[12]), .B(arg[15]), .C(n946), .D(n945), .Q(n947) );
  INV6 U1306 ( .A(n1287), .Q(n1300) );
  NOR33 U1307 ( .A(n1224), .B(n1142), .C(n1141), .Q(n903) );
  INV6 U1308 ( .A(n1127), .Q(n1115) );
  INV15 U1309 ( .A(arg[14]), .Q(n925) );
  OAI212 U1310 ( .A(n1390), .B(n1389), .C(n767), .Q(n1391) );
  OAI312 U1311 ( .A(n1336), .B(n1335), .C(n1334), .D(n1333), .Q(n1354) );
  NAND22 U1312 ( .A(n1274), .B(n1278), .Q(n1301) );
  NAND22 U1313 ( .A(arg[2]), .B(n858), .Q(n859) );
  INV3 U1314 ( .A(n1253), .Q(n858) );
  OAI211 U1315 ( .A(n888), .B(n1248), .C(lt_gt_52_A_1_), .Q(n1253) );
  OAI2111 U1316 ( .A(n716), .B(n888), .C(n1430), .D(n1340), .Q(n1252) );
  OAI212 U1317 ( .A(n1364), .B(n699), .C(n1363), .Q(n1451) );
  INV15 U1318 ( .A(n886), .Q(lt_gt_52_A_4_) );
  INV0 U1319 ( .A(n727), .Q(n1357) );
  AOI212 U1320 ( .A(n1396), .B(n878), .C(n1452), .Q(n1397) );
  OAI222 U1321 ( .A(n1416), .B(n1415), .C(n1416), .D(n1414), .Q(n1417) );
  OAI212 U1322 ( .A(lt_gt_52_A_4_), .B(n1395), .C(n1446), .Q(n1447) );
  OAI222 U1323 ( .A(n1266), .B(n1265), .C(n878), .D(n1353), .Q(n1267) );
  NAND22 U1324 ( .A(n862), .B(N718), .Q(n1468) );
  IMUX24 U1325 ( .A(n904), .B(n1223), .S(lt_gt_52_A_1_), .Q(n1350) );
  NAND24 U1326 ( .A(n1234), .B(n1210), .Q(n1269) );
  IMUX24 U1327 ( .A(n1171), .B(n1170), .S(n1169), .Q(n1286) );
  OAI212 U1328 ( .A(n1133), .B(n827), .C(n668), .Q(n1281) );
  NAND20 U1329 ( .A(n1406), .B(n879), .Q(n1407) );
  OAI212 U1330 ( .A(n878), .B(n1353), .C(n1242), .Q(n1243) );
  CLKIN1 U1331 ( .A(n865), .Q(n965) );
  AOI312 U1332 ( .A(n1018), .B(n1003), .C(n1058), .D(n1002), .Q(n863) );
  NAND28 U1333 ( .A(n981), .B(n864), .Q(n944) );
  NAND28 U1334 ( .A(n814), .B(arg[14]), .Q(n955) );
  INV15 U1335 ( .A(arg[14]), .Q(n930) );
  INV4 U1336 ( .A(n1312), .Q(n1316) );
  AOI312 U1337 ( .A(n1198), .B(n1197), .C(n1196), .D(n1195), .Q(n1199) );
  NAND21 U1338 ( .A(n1459), .B(n1458), .Q(n1449) );
  AOI2112 U1339 ( .A(roundup), .B(n1460), .C(n1461), .D(n1455), .Q(n1456) );
  CLKIN0 U1340 ( .A(n755), .Q(n1165) );
  AOI210 U1341 ( .A(n1358), .B(n908), .C(n1357), .Q(n1368) );
  INV3 U1342 ( .A(n1461), .Q(n1462) );
  INV3 U1343 ( .A(n873), .Q(lt_gt_52_A_7_) );
  CLKIN3 U1344 ( .A(arg[12]), .Q(n870) );
  OAI212 U1345 ( .A(n998), .B(n997), .C(n920), .Q(n999) );
  XNR20 U1346 ( .A(lt_gt_52_A_1_), .B(n1430), .Q(n1433) );
  INV3 U1347 ( .A(arg[4]), .Q(n1206) );
  NOR20 U1348 ( .A(n1470), .B(n1433), .Q(n874) );
  INV3 U1349 ( .A(n874), .Q(n875) );
  CLKIN2 U1350 ( .A(N711), .Q(n894) );
  CLKIN2 U1351 ( .A(N716), .Q(n900) );
  INV3 U1352 ( .A(n1123), .Q(n1137) );
  INV3 U1353 ( .A(n1083), .Q(n1086) );
  INV3 U1354 ( .A(n1435), .Q(n1429) );
  XNR21 U1355 ( .A(n1122), .B(n1121), .Q(n877) );
  INV3 U1356 ( .A(arg[5]), .Q(n1210) );
  XNR22 U1357 ( .A(arg[10]), .B(n949), .Q(n989) );
  INV3 U1358 ( .A(N712), .Q(n897) );
  INV3 U1359 ( .A(N715), .Q(n899) );
  NAND22 U1360 ( .A(n1177), .B(n1202), .Q(n1184) );
  MUX21 U1361 ( .A(N713), .B(n888), .S(n1466), .Q(sqroot[3]) );
  MUX21 U1362 ( .A(N714), .B(lt_gt_52_A_4_), .S(n1466), .Q(sqroot[4]) );
  MUX21 U1363 ( .A(N717), .B(n908), .S(n1466), .Q(sqroot[7]) );
  BUF2 U1364 ( .A(lt_gt_52_A_7_), .Q(n908) );
  AOI220 U1365 ( .A(n887), .B(n1081), .C(n1080), .D(n1079), .Q(n1089) );
  AOI220 U1366 ( .A(n887), .B(n1087), .C(n1086), .D(n1085), .Q(n1088) );
  NOR20 U1367 ( .A(n1224), .B(n831), .Q(n1227) );
  AOI210 U1368 ( .A(n1209), .B(n1206), .C(n888), .Q(n1208) );
  NAND21 U1369 ( .A(arg[11]), .B(n962), .Q(n967) );
  NAND22 U1370 ( .A(n963), .B(arg[11]), .Q(n956) );
  LOGIC0 U1371 ( .Q(n1472) );
  NAND34 U1372 ( .A(n1120), .B(n1119), .C(n1122), .Q(n1109) );
  NAND33 U1373 ( .A(n1180), .B(n1156), .C(n1155), .Q(n1177) );
  OAI212 U1374 ( .A(n737), .B(n1401), .C(n1400), .Q(n1465) );
  AOI311 U1375 ( .A(n869), .B(n1362), .C(n1385), .D(n1360), .Q(n1363) );
  AOI2112 U1376 ( .A(n1322), .B(n1172), .C(n1273), .D(n911), .Q(n1204) );
  NAND43 U1377 ( .A(n1087), .B(n1137), .C(n1110), .D(n1109), .Q(n892) );
  INV1 U1378 ( .A(n1468), .Q(sqroot[8]) );
  NAND32 U1379 ( .A(n1119), .B(n863), .C(n706), .Q(n1073) );
  OAI222 U1380 ( .A(n1189), .B(n1095), .C(n1094), .D(n1093), .Q(n893) );
  OAI2112 U1381 ( .A(n728), .B(n802), .C(n1096), .D(n1090), .Q(n1094) );
  IMUX20 U1382 ( .A(n894), .B(n895), .S(n1466), .Q(sqroot[1]) );
  IMUX20 U1383 ( .A(n897), .B(n898), .S(n1466), .Q(sqroot[2]) );
  IMUX20 U1384 ( .A(n899), .B(n909), .S(n1466), .Q(sqroot[5]) );
  IMUX20 U1385 ( .A(n900), .B(n694), .S(n1466), .Q(sqroot[6]) );
  NAND28 U1386 ( .A(n1092), .B(n1091), .Q(n1179) );
  AOI2111 U1387 ( .A(n1176), .B(n1197), .C(n1195), .D(n1175), .Q(n1187) );
  BUF2 U1388 ( .A(n695), .Q(n904) );
  XNR20 U1389 ( .A(n902), .B(arg[7]), .Q(n1118) );
  IMUX24 U1390 ( .A(n1165), .B(n1164), .S(n1169), .Q(n1285) );
  INV6 U1391 ( .A(n1280), .Q(n1284) );
  IMUX24 U1392 ( .A(n1227), .B(n1226), .S(n1240), .Q(n1405) );
  OAI211 U1393 ( .A(n932), .B(n931), .C(n1403), .Q(n935) );
  NAND28 U1394 ( .A(n680), .B(n1244), .Q(n1228) );
  NAND26 U1395 ( .A(n917), .B(n916), .Q(n964) );
  NOR41 U1396 ( .A(n1271), .B(n1270), .C(n1273), .D(n1269), .Q(n1272) );
  NOR42 U1397 ( .A(n1450), .B(n1337), .C(n1454), .D(n1356), .Q(n1349) );
  INV6 U1398 ( .A(n1305), .Q(n1335) );
  NOR33 U1399 ( .A(n1066), .B(n1105), .C(n1104), .Q(n1067) );
  NOR42 U1400 ( .A(n741), .B(n854), .C(n932), .D(n931), .Q(n958) );
  INV6 U1401 ( .A(n929), .Q(n931) );
  NOR42 U1402 ( .A(n1450), .B(n1101), .C(n1010), .D(n1001), .Q(n1002) );
  NAND43 U1403 ( .A(n1012), .B(n988), .C(n987), .D(n756), .Q(n1021) );
  OAI222 U1404 ( .A(n644), .B(n856), .C(arg[13]), .D(arg[15]), .Q(n915) );
  CLKIN3 U1405 ( .A(arg[9]), .Q(n918) );
  OAI312 U1406 ( .A(arg[14]), .B(arg[12]), .C(arg[13]), .D(n955), .Q(n1403) );
  OAI212 U1407 ( .A(arg[11]), .B(n991), .C(n911), .Q(n996) );
  AOI212 U1408 ( .A(n1008), .B(n910), .C(n920), .Q(n923) );
  OAI212 U1409 ( .A(n909), .B(n1008), .C(n921), .Q(n922) );
  OAI222 U1410 ( .A(arg[14]), .B(n945), .C(arg[12]), .D(arg[15]), .Q(n952) );
  CLKIN3 U1411 ( .A(n952), .Q(n936) );
  AOI312 U1412 ( .A(arg[13]), .B(n927), .C(n926), .D(n944), .Q(n932) );
  OAI212 U1413 ( .A(arg[15]), .B(n930), .C(arg[12]), .Q(n928) );
  OAI2112 U1414 ( .A(arg[13]), .B(arg[14]), .C(n928), .D(n944), .Q(n929) );
  OAI212 U1415 ( .A(arg[11]), .B(n909), .C(n938), .Q(n939) );
  OAI212 U1416 ( .A(arg[12]), .B(n941), .C(arg[13]), .Q(n942) );
  OAI312 U1417 ( .A(n741), .B(n943), .C(n1172), .D(n942), .Q(n948) );
  OAI212 U1418 ( .A(arg[14]), .B(arg[15]), .C(n944), .Q(n946) );
  OAI2112 U1419 ( .A(n952), .B(n953), .C(n954), .D(lt_gt_52_A_7_), .Q(n1006)
         );
  OAI212 U1420 ( .A(arg[12]), .B(arg[13]), .C(n955), .Q(n962) );
  OAI212 U1421 ( .A(n961), .B(n960), .C(n959), .Q(n969) );
  AOI2112 U1422 ( .A(n964), .B(n965), .C(arg[10]), .D(n963), .Q(n966) );
  NOR33 U1423 ( .A(n970), .B(n968), .C(n969), .Q(n1007) );
  OAI212 U1424 ( .A(n974), .B(n973), .C(n972), .Q(n975) );
  CLKIN3 U1425 ( .A(n1008), .Q(n982) );
  OAI212 U1426 ( .A(n991), .B(n911), .C(n985), .Q(n983) );
  NAND22 U1427 ( .A(n911), .B(n1008), .Q(n984) );
  OAI312 U1428 ( .A(n911), .B(n997), .C(n998), .D(n891), .Q(n1009) );
  AOI2112 U1429 ( .A(n994), .B(n1450), .C(n911), .D(n993), .Q(n1003) );
  AOI312 U1430 ( .A(n711), .B(n1004), .C(n1003), .D(n1002), .Q(n1107) );
  OAI212 U1431 ( .A(n1008), .B(n1026), .C(n1025), .Q(n1033) );
  OAI212 U1432 ( .A(n692), .B(n1011), .C(n736), .Q(n1014) );
  AOI212 U1433 ( .A(n1014), .B(n1450), .C(n1064), .Q(n1015) );
  CLKIN3 U1434 ( .A(arg[6]), .Q(n1122) );
  NAND22 U1435 ( .A(n1087), .B(n1122), .Q(n1081) );
  CLKIN3 U1436 ( .A(n1081), .Q(n1035) );
  OAI2112 U1437 ( .A(n908), .B(n710), .C(n1019), .D(n1020), .Q(n1063) );
  NAND22 U1438 ( .A(n1025), .B(n1035), .Q(n1030) );
  OAI212 U1439 ( .A(n1072), .B(n1061), .C(n1039), .Q(n1075) );
  OAI2112 U1440 ( .A(n1061), .B(n1072), .C(n1039), .D(n879), .Q(n1040) );
  OAI312 U1441 ( .A(n911), .B(n1043), .C(n1042), .D(n1041), .Q(n1044) );
  AOI312 U1442 ( .A(n1046), .B(n823), .C(n705), .D(n1045), .Q(n1047) );
  OAI212 U1443 ( .A(n802), .B(n1053), .C(n1052), .Q(n1054) );
  NAND22 U1444 ( .A(n1179), .B(n908), .Q(n1095) );
  CLKIN3 U1445 ( .A(n1078), .Q(n1084) );
  OAI212 U1446 ( .A(arg[6]), .B(n1087), .C(n1084), .Q(n1080) );
  NAND22 U1447 ( .A(n1210), .B(n1206), .Q(n1123) );
  NAND22 U1448 ( .A(n1137), .B(n1122), .Q(n1083) );
  NAND22 U1449 ( .A(n1083), .B(n1122), .Q(n1079) );
  NAND22 U1450 ( .A(arg[7]), .B(n1084), .Q(n1085) );
  OAI222 U1451 ( .A(n1189), .B(n1095), .C(n1093), .D(n688), .Q(n1130) );
  OAI212 U1452 ( .A(n908), .B(n1179), .C(n1096), .Q(n1127) );
  OAI222 U1453 ( .A(n1171), .B(n823), .C(n1097), .D(n746), .Q(n1099) );
  OAI2112 U1454 ( .A(arg[6]), .B(n1137), .C(n1124), .D(n1057), .Q(n1152) );
  OAI222 U1455 ( .A(n1138), .B(n1206), .C(n893), .D(n1129), .Q(n1131) );
  CLKIN3 U1456 ( .A(arg[3]), .Q(n1257) );
  CLKIN3 U1457 ( .A(arg[2]), .Q(n1340) );
  NAND22 U1458 ( .A(n1257), .B(n1340), .Q(n1235) );
  AOI2112 U1459 ( .A(n1132), .B(arg[4]), .C(n1235), .D(n1131), .Q(n1234) );
  CLKIN3 U1460 ( .A(n1235), .Q(n1209) );
  OAI2112 U1461 ( .A(arg[4]), .B(n1209), .C(n1140), .D(n1470), .Q(n1237) );
  OAI222 U1462 ( .A(n1145), .B(n1225), .C(n903), .D(n888), .Q(n1274) );
  OAI212 U1463 ( .A(n687), .B(n754), .C(n1177), .Q(n1173) );
  OAI312 U1464 ( .A(n737), .B(n722), .C(n1153), .D(n1152), .Q(n1167) );
  AOI212 U1465 ( .A(n1158), .B(n1197), .C(n1175), .Q(n1162) );
  CLKIN3 U1466 ( .A(n1307), .Q(n1191) );
  OAI222 U1467 ( .A(n1308), .B(n1307), .C(n1191), .D(n1190), .Q(n1192) );
  CLKIN3 U1468 ( .A(n1218), .Q(n1295) );
  NOR24 U1469 ( .A(n1295), .B(n1296), .Q(n1203) );
  OAI2112 U1470 ( .A(n696), .B(n1204), .C(n1203), .D(n1332), .Q(n1205) );
  OAI312 U1471 ( .A(n1208), .B(n1224), .C(n831), .D(n1216), .Q(n1214) );
  AOI2112 U1472 ( .A(n901), .B(n887), .C(n1213), .D(n1214), .Q(n1215) );
  OAI222 U1473 ( .A(n878), .B(n1286), .C(n908), .D(n1285), .Q(n1220) );
  AOI2112 U1474 ( .A(n668), .B(n910), .C(n1219), .D(n1220), .Q(n1221) );
  AOI312 U1475 ( .A(lt_gt_52_A_4_), .B(n1231), .C(n700), .D(n1229), .Q(n1232)
         );
  CLKIN3 U1476 ( .A(arg[1]), .Q(n1250) );
  CLKIN3 U1477 ( .A(arg[0]), .Q(n1249) );
  NAND22 U1478 ( .A(n1250), .B(n1249), .Q(n1251) );
  CLKIN3 U1479 ( .A(n1251), .Q(n1430) );
  OAI212 U1480 ( .A(n888), .B(n716), .C(n1384), .Q(n1261) );
  AOI212 U1481 ( .A(n1277), .B(n1302), .C(n1276), .Q(n1279) );
  NAND22 U1482 ( .A(n1291), .B(n910), .Q(n1312) );
  OAI212 U1483 ( .A(n909), .B(n768), .C(n1314), .Q(n1330) );
  OAI2112 U1484 ( .A(n1450), .B(n1292), .C(n746), .D(n1317), .Q(n1305) );
  AOI312 U1485 ( .A(n1329), .B(n1305), .C(n1304), .D(n1331), .Q(n1306) );
  OAI212 U1486 ( .A(n895), .B(n1310), .C(n1309), .Q(n1369) );
  OAI212 U1487 ( .A(n1316), .B(n1315), .C(n1314), .Q(n1320) );
  AOI212 U1488 ( .A(n1320), .B(n1319), .C(n1318), .Q(n1321) );
  OAI312 U1489 ( .A(n1325), .B(n852), .C(n1324), .D(n1323), .Q(n1356) );
  AOI2112 U1490 ( .A(n1454), .B(n1450), .C(n1369), .D(n727), .Q(n1326) );
  OAI212 U1491 ( .A(n1328), .B(n1327), .C(n1326), .Q(n1373) );
  OAI222 U1492 ( .A(arg[2]), .B(n1430), .C(lt_gt_52_A_1_), .D(n1340), .Q(n1410) );
  AOI312 U1493 ( .A(n1388), .B(n685), .C(n1342), .D(n634), .Q(n1344) );
  OAI212 U1494 ( .A(n1346), .B(n1345), .C(n699), .Q(n1348) );
  OAI212 U1495 ( .A(n1375), .B(n767), .C(n1374), .Q(n1376) );
  CLKIN3 U1496 ( .A(roundup), .Q(n1452) );
  AOI312 U1497 ( .A(n1427), .B(n1428), .C(n1426), .D(n1425), .Q(n1439) );
  NAND24 U1498 ( .A(n1429), .B(n898), .Q(n1432) );
  OAI222 U1499 ( .A(n1439), .B(n1438), .C(n1436), .D(n898), .Q(n1440) );
  XNR21 U1500 ( .A(n1451), .B(n1450), .Q(n1453) );
  OAI2112 U1501 ( .A(n1465), .B(n1464), .C(n1463), .D(n1462), .Q(n1467) );
endmodule

